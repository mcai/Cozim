// $Id: vcr_sw_alloc_sep_if.v 5188 2012-08-30 00:31:31Z dub $

/*
 Copyright (c) 2007-2012, Trustees of The Leland Stanford Junior University
 All rights reserved.

 Redistribution and use in source and binary forms, with or without
 modification, are permitted provided that the following conditions are met:

 Redistributions of source code must retain the above copyright notice, this 
 list of conditions and the following disclaimer.
 Redistributions in binary form must reproduce the above copyright notice, this
 list of conditions and the following disclaimer in the documentation and/or
 other materials provided with the distribution.

 THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
 ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
 WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE 
 DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR
 ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
 (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
 LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON
 ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
 (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
 SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/

//==============================================================================
// switch allocator variant using separable input-first allocation
//==============================================================================

module vcr_sw_alloc_sep_if
  (clk, reset, active_ip, active_op, route_ip_ivc_op, req_nonspec_ip_ivc, 
   req_spec_ip_ivc, gnt_ip, sel_ip_ivc, gnt_op, sel_op_ip, sel_op_ivc);
   
`include "clib/c_functions.sv"
`include "clib/c_constants.sv"
`include "vcr_constants.sv"
   
   // number of VCs
   parameter num_vcs = 4;
   
   // number of input and output ports on switch
   parameter num_ports = 5;
   
   // select which arbiter type to use in allocator
   parameter arbiter_type = `ARBITER_TYPE_ROUND_ROBIN_BINARY;
   
   // select speculation type
   parameter spec_type = `SW_ALLOC_SPEC_TYPE_REQ;
   
   parameter reset_type = `RESET_TYPE_ASYNC;
   
   input clk;
   input reset;
   
   // clock enable signals
   input [0:num_ports-1] active_ip;
   input [0:num_ports-1] active_op;
   
   // destination port selects
   input [0:num_ports*num_vcs*num_ports-1] route_ip_ivc_op;
   
   // non-speculative switch requests
   input [0:num_ports*num_vcs-1] 	   req_nonspec_ip_ivc;
   
   // speculative switch requests
   input [0:num_ports*num_vcs-1] 	   req_spec_ip_ivc;
   
   // grants
   output [0:num_ports-1] 		   gnt_ip;
   wire [0:num_ports-1] 		   gnt_ip;
   
   // indicate which VC at a given port is granted
   output [0:num_ports*num_vcs-1] 	   sel_ip_ivc;
   wire [0:num_ports*num_vcs-1] 	   sel_ip_ivc;
   
   // grants for output ports
   output [0:num_ports-1] 		   gnt_op;
   wire [0:num_ports-1] 		   gnt_op;
   
   // selected input ports (if any)
   output [0:num_ports*num_ports-1] 	   sel_op_ip;
   wire [0:num_ports*num_ports-1] 	   sel_op_ip;
   
   // selected input VCs (if any)
   output [0:num_ports*num_vcs-1] 	   sel_op_ivc;
   wire [0:num_ports*num_vcs-1] 	   sel_op_ivc;
   
   
   //---------------------------------------------------------------------------
   // global wires
   //---------------------------------------------------------------------------
   
   wire [0:num_ports*num_ports-1] 	   req_in_nonspec_ip_op;   
   wire [0:num_ports*num_ports-1] 	   req_out_nonspec_ip_op;
   wire [0:num_ports*num_ports-1] 	   gnt_out_nonspec_ip_op;
   
   wire [0:num_ports*num_ports-1] 	   req_out_spec_ip_op;
   wire [0:num_ports*num_ports-1] 	   gnt_out_spec_ip_op;
   
   wire [0:num_ports-1] 		   unused_by_nonspec_ip;
   wire [0:num_ports-1] 		   unused_by_nonspec_op;
   
   
   //---------------------------------------------------------------------------
   // input stage
   //---------------------------------------------------------------------------
   
   generate
      
      genvar 				   ip;
      
      for(ip = 0; ip < num_ports; ip = ip + 1)
	begin:ips
	   
	   wire active;
	   assign active = active_ip[ip];
	   
	   wire [0:num_vcs*num_ports-1] route_ivc_op;
	   assign route_ivc_op
	     = route_ip_ivc_op[ip*num_vcs*num_ports:(ip+1)*num_vcs*num_ports-1];
	   
	   
	   //-------------------------------------------------------------------
	   // perform input-side arbitration
	   //-------------------------------------------------------------------
	   
	   wire [0:num_ports-1] 	gnt_out_nonspec_op;
	   assign gnt_out_nonspec_op
	     = gnt_out_nonspec_ip_op[ip*num_ports:(ip+1)*num_ports-1];
	   
	   wire 			gnt_out_nonspec;
	   assign gnt_out_nonspec = |gnt_out_nonspec_op;
	   
	   wire 			update_arb_nonspec;
	   assign update_arb_nonspec = gnt_out_nonspec;
	   
	   wire [0:num_vcs-1] 		req_nonspec_ivc;
	   assign req_nonspec_ivc
	     = req_nonspec_ip_ivc[ip*num_vcs:(ip+1)*num_vcs-1];
	   
	   wire [0:num_vcs-1] 		req_in_nonspec_ivc;
	   assign req_in_nonspec_ivc = req_nonspec_ivc;
	   
	   wire [0:num_vcs-1] 		gnt_in_nonspec_ivc;
	   
	   if(spec_type != `SW_ALLOC_SPEC_TYPE_PRIO)
	     begin
		
		c_arbiter
		  #(.num_ports(num_vcs),
		    .num_priorities(1),
		    .reset_type(reset_type),
		    .arbiter_type(arbiter_type))
		gnt_in_nonspec_ivc_arb
		  (.clk(clk),
		   .reset(reset),
		   .active(active),
		   .update(update_arb_nonspec),
		   .req_pr(req_in_nonspec_ivc),
		   .gnt_pr(gnt_in_nonspec_ivc),
		   .gnt());
		
	     end
	   
	   wire [0:num_ports-1] req_in_nonspec_op;
	   c_select_mofn
	     #(.width(num_ports),
	       .num_ports(num_vcs))
	   req_in_nonspec_ip_op_sel
	     (.select(req_in_nonspec_ivc),
	      .data_in(route_ivc_op),
	      .data_out(req_in_nonspec_op));
	   
	   assign req_in_nonspec_ip_op[ip*num_ports:(ip+1)*num_ports-1]
	     = req_in_nonspec_op;
	   
	   //-------------------------------------------------------------------
	   // generate requests for output stage
	   //-------------------------------------------------------------------
	   
	   wire [0:num_ports-1] req_out_nonspec_op;
	   c_select_mofn
	     #(.width(num_ports),
	       .num_ports(num_vcs))
	   req_out_nonspec_op_sel
	     (.select(gnt_in_nonspec_ivc),
	      .data_in(route_ivc_op),
	      .data_out(req_out_nonspec_op));
	   
	   assign req_out_nonspec_ip_op[ip*num_ports:(ip+1)*num_ports-1]
	     = req_out_nonspec_op;
	   
	   
	   //-------------------------------------------------------------------
	   // handle speculative requests
	   //-------------------------------------------------------------------
	   
	   wire [0:num_ports-1] req_out_spec_op;
	   wire 		gnt;
	   wire [0:num_vcs-1] 	sel_ivc;
	   
	   if(spec_type != `SW_ALLOC_SPEC_TYPE_NONE)
	     begin
		
		//--------------------------------------------------------------
		// perform input-side arbitration (speculative)
		//--------------------------------------------------------------
		
		wire [0:num_ports-1] gnt_out_spec_op;
		assign gnt_out_spec_op
		  = gnt_out_spec_ip_op[ip*num_ports:(ip+1)*num_ports-1];
		
		wire 		     gnt_out_spec;
		assign gnt_out_spec = |gnt_out_spec_op;
		
		wire 		     update_arb_spec;
		assign update_arb_spec = gnt_out_spec;
		
		wire [0:num_vcs-1]   req_spec_ivc;
		assign req_spec_ivc
		  = req_spec_ip_ivc[ip*num_vcs:(ip+1)*num_vcs-1];
		
		wire [0:num_vcs-1]   req_in_spec_ivc;
		assign req_in_spec_ivc = req_spec_ivc;
		
		wire [0:num_vcs-1]   gnt_in_spec_ivc;
		
		if(spec_type == `SW_ALLOC_SPEC_TYPE_PRIO)
		  begin
		     
		     wire update_arb;
		     assign update_arb = update_arb_spec | update_arb_nonspec;
		     
		     c_arbiter
		       #(.num_ports(num_vcs),
			 .num_priorities(2),
			 .reset_type(reset_type),
			 .arbiter_type(arbiter_type))
		     gnt_in_ivc_arb
		       (.clk(clk),
			.reset(reset),
			.active(active),
			.update(update_arb),
			.req_pr({req_in_nonspec_ivc, req_in_spec_ivc}),
			.gnt_pr({gnt_in_nonspec_ivc, gnt_in_spec_ivc}),
			.gnt(sel_ivc));
		     
		     assign gnt = gnt_out_nonspec | gnt_out_spec;
		     
		  end
		else
		  begin
		     
		     c_arbiter
		       #(.num_ports(num_vcs),
			 .num_priorities(1),
			 .reset_type(reset_type),
			 .arbiter_type(arbiter_type))
		     gnt_in_spec_ivc_arb
		       (.clk(clk),
			.reset(reset),
			.active(active),
			.update(update_arb_spec),
			.req_pr(req_in_spec_ivc),
			.gnt_pr(gnt_in_spec_ivc),
			.gnt());
		     
		     wire unused_by_nonspec;
		     assign unused_by_nonspec = unused_by_nonspec_ip[ip];
		     
		     wire [0:num_ports-1] gnt_out_spec_qual_op;
		     assign gnt_out_spec_qual_op
		       = gnt_out_spec_op & unused_by_nonspec_op &
			 {num_ports{unused_by_nonspec}};
		     
		     wire 		  gnt_out_spec_qual;
		     assign gnt_out_spec_qual = |gnt_out_spec_qual_op;
		     
		     assign gnt = gnt_out_nonspec | gnt_out_spec_qual;
		     
		     case(spec_type)
		       
		       `SW_ALLOC_SPEC_TYPE_REQ:
			 begin
			    
			    wire req_nonspec;
			    assign req_nonspec = |req_nonspec_ivc;
			    
			    assign sel_ivc = req_nonspec ? 
					     gnt_in_nonspec_ivc : 
					     gnt_in_spec_ivc;
			    
			 end
		       
		       `SW_ALLOC_SPEC_TYPE_GNT:
			 begin
			    
			    assign sel_ivc = gnt_out_nonspec ? 
					     gnt_in_nonspec_ivc : 
					     gnt_in_spec_ivc;
			    
			 end
		       
		     endcase
		     
		  end
		
		
		//--------------------------------------------------------------
		// generate requests for output stage (speculative)
		//--------------------------------------------------------------
		
		c_select_mofn
		  #(.width(num_ports),
		    .num_ports(num_vcs))
		req_out_spec_op_sel
		  (.select(gnt_in_spec_ivc),
		   .data_in(route_ivc_op),
		   .data_out(req_out_spec_op));
		
	     end
	   else
	     begin
		
		assign req_out_spec_op = {num_ports{1'b0}};
		assign sel_ivc = gnt_in_nonspec_ivc;
		assign gnt = gnt_out_nonspec;
		
	     end
	   
	   
	   //-------------------------------------------------------------------
	   // combine global grants
	   //-------------------------------------------------------------------
	   
	   assign req_out_spec_ip_op[ip*num_ports:(ip+1)*num_ports-1]
	     = req_out_spec_op;
	   assign sel_ip_ivc[ip*num_vcs:(ip+1)*num_vcs-1] = sel_ivc;
	   assign gnt_ip[ip] = gnt;
	   	   
	end
      
   endgenerate
   
   
   //---------------------------------------------------------------------------
   // bit shuffling for changing sort order
   //---------------------------------------------------------------------------
   
   wire [0:num_ports*num_ports-1] req_in_nonspec_op_ip;
   c_interleave
     #(.width(num_ports*num_ports),
       .num_blocks(num_ports))
   req_in_nonspec_op_ip_intl
     (.data_in(req_in_nonspec_ip_op),
      .data_out(req_in_nonspec_op_ip));
   
   wire [0:num_ports*num_ports-1] req_out_nonspec_op_ip;
   c_interleave
     #(.width(num_ports*num_ports),
       .num_blocks(num_ports))
   req_out_nonspec_op_ip_intl
     (.data_in(req_out_nonspec_ip_op),
      .data_out(req_out_nonspec_op_ip));
   
   wire [0:num_ports*num_ports-1] gnt_out_nonspec_op_ip;
   c_interleave
     #(.width(num_ports*num_ports),
       .num_blocks(num_ports))
   gnt_out_nonspec_op_ip_intl
     (.data_in(gnt_out_nonspec_op_ip),
      .data_out(gnt_out_nonspec_ip_op));
   
   wire [0:num_ports*num_ports-1] req_out_spec_op_ip;
   c_interleave
     #(.width(num_ports*num_ports),
       .num_blocks(num_ports))
   req_out_spec_op_ip_intl
     (.data_in(req_out_spec_ip_op),
      .data_out(req_out_spec_op_ip));
   
   wire [0:num_ports*num_ports-1] gnt_out_spec_op_ip;
   c_interleave
     #(.width(num_ports*num_ports),
       .num_blocks(num_ports))
   gnt_out_spec_op_ip_intl
     (.data_in(gnt_out_spec_op_ip),
      .data_out(gnt_out_spec_ip_op));
   
   
   //---------------------------------------------------------------------------
   // mask speculative requests that conflict with non-speculative ones
   //---------------------------------------------------------------------------
   
   generate
      
      case(spec_type)
	
	`SW_ALLOC_SPEC_TYPE_NONE, `SW_ALLOC_SPEC_TYPE_PRIO:
	  begin
	     
	     assign unused_by_nonspec_ip = {num_ports{1'b0}};
	     assign unused_by_nonspec_op = {num_ports{1'b0}};
	     
	  end
	
	`SW_ALLOC_SPEC_TYPE_REQ:
	  begin
	     
	     // We can potentially improve matching by using the grants of the
	     // input stage (i.e., the requests of the output stage) to filter 
	     // out output ports that have all requests for them eliminated in 
	     // the input stage. As the associated OR reduction can be performed
	     // in parallel with output-stage arbitration, this should not 
	     // increase delay.
	     c_binary_op
	       #(.width(num_ports),
		 .num_ports(num_ports),
		 .op(`BINARY_OP_NOR))
	     unused_by_nonspec_op_nor
	       (.data_in(req_out_nonspec_ip_op),
		.data_out(unused_by_nonspec_op));
	     
	     // For determining which inputs are in use, looking at the input-
	     // stage grants rather than its requests does not yield any 
	     // additional information, as the input-side arbitration stage will
	     // generate a grant if and only if there were any requests. Thus,
	     // we use the requests here to ease timing.
	     c_binary_op
	       #(.width(num_ports),
		 .num_ports(num_ports),
		 .op(`BINARY_OP_NOR))
	     unused_by_nonspec_ip_nor
	       (.data_in(req_in_nonspec_op_ip),
		.data_out(unused_by_nonspec_ip));
	     
	  end
	
	`SW_ALLOC_SPEC_TYPE_GNT:
	  begin
	     
	     // An output is granted if and only if there were any output-stage 
	     // requests for it; thus, it is sufficient to look at the arbiter 
	     // inputs here.
	     c_binary_op
	       #(.width(num_ports),
		 .num_ports(num_ports),
		 .op(`BINARY_OP_NOR))
	     unused_by_nonspec_op_nor
	       (.data_in(req_out_nonspec_ip_op),
		.data_out(unused_by_nonspec_op));
	     
	     // However, we can make no such simplification to determine which
	     // input ports are in use: A given input may have requested 
	     // one or more outputs, but all of its requests could have been 
	     // eliminated in the output arbitration stage.
	     c_binary_op
	       #(.width(num_ports),
		 .num_ports(num_ports),
		 .op(`BINARY_OP_NOR))
	     unused_by_nonspec_ip_nor
	       (.data_in(gnt_out_nonspec_op_ip),
		.data_out(unused_by_nonspec_ip));
	     
	  end
	
      endcase
      
   endgenerate
   
   
   //---------------------------------------------------------------------------
   // output stage
   //---------------------------------------------------------------------------
   
   generate
      
      genvar 				    op;
      
      for (op = 0; op < num_ports; op = op + 1)
	begin:ops
	   
	   wire active;
	   assign active = active_op[op];
	   
	   
	   //-------------------------------------------------------------------
	   // perform output-side arbitration (select input port)
	   //-------------------------------------------------------------------
	   
	   wire [0:num_ports-1] sel_ip;
	   
	   wire [0:num_ports-1] req_out_nonspec_ip;
	   assign req_out_nonspec_ip
	     = req_out_nonspec_op_ip[op*num_ports:(op+1)*num_ports-1];
	   
	   wire req_out_nonspec;
	   assign req_out_nonspec = |req_out_nonspec_ip;
	   
	   // if any VC requesting this output port was granted at any input
	   // port in the first stage, one of these input ports will be granted
	   // here as well, and we can thus update priorities
	   wire 		update_arb_nonspec;
	   assign update_arb_nonspec = req_out_nonspec;
	   
	   wire [0:num_ports-1] gnt_out_nonspec_ip;
	   
	   if(spec_type != `SW_ALLOC_SPEC_TYPE_PRIO)
	     begin
		
		c_arbiter
		  #(.num_ports(num_ports),
		    .num_priorities(1),
		    .arbiter_type(arbiter_type),
		    .reset_type(reset_type))
		gnt_out_nonspec_ip_arb
		  (.clk(clk),
		   .reset(reset),
		   .active(active),
		   .update(update_arb_nonspec),
		   .req_pr(req_out_nonspec_ip),
		   .gnt_pr(gnt_out_nonspec_ip),
		   .gnt());
		
	     end
	   
	   
	   //-------------------------------------------------------------------
	   // handle speculative requests
	   //-------------------------------------------------------------------
	   
	   wire [0:num_ports-1] gnt_out_spec_ip;
	   wire 		gnt;
	   
	   if(spec_type != `SW_ALLOC_SPEC_TYPE_NONE)
	     begin
		
		//--------------------------------------------------------------
		// perform output-side arbitration (speculative)
		//--------------------------------------------------------------
		
		wire [0:num_ports-1] req_out_spec_ip;
		assign req_out_spec_ip
		  = req_out_spec_op_ip[op*num_ports:(op+1)*num_ports-1];

		wire 		     req_out_spec;
		assign req_out_spec = |req_out_spec_ip;
		
		wire 		     update_arb_spec;
		assign update_arb_spec = req_out_spec;
		
		if(spec_type == `SW_ALLOC_SPEC_TYPE_PRIO)
		  begin
		     
		     wire update_arb;
		     assign update_arb = update_arb_nonspec | update_arb_spec;
		     
		     c_arbiter
		       #(.num_ports(num_ports),
			 .num_priorities(2),
			 .arbiter_type(arbiter_type),
			 .reset_type(reset_type))
		     gnt_out_ip_arb
		       (.clk(clk),
			.reset(reset),
			.active(active),
			.update(update_arb),
			.req_pr({req_out_nonspec_ip, req_out_spec_ip}),
			.gnt_pr({gnt_out_nonspec_ip, gnt_out_spec_ip}),
			.gnt(sel_ip));
		     
		     assign gnt = req_out_nonspec | req_out_spec;
		     
		  end
		else
		  begin
		     
		     c_arbiter
		       #(.num_ports(num_ports),
			 .num_priorities(1),
			 .arbiter_type(arbiter_type),
			 .reset_type(reset_type))
		     gnt_out_spec_ip_arb
		       (.clk(clk),
			.reset(reset),
			.active(active),
			.update(update_arb_spec),
			.req_pr(req_out_spec_ip),
			.gnt_pr(gnt_out_spec_ip),
			.gnt());
		     
		     wire unused_by_nonspec;
		     assign unused_by_nonspec = unused_by_nonspec_op[op];
		     
		     wire [0:num_ports-1] gnt_out_spec_qual_ip;
		     assign gnt_out_spec_qual_ip
		       = gnt_out_spec_ip & unused_by_nonspec_ip &
			 {num_ports{unused_by_nonspec}};
		     
		     wire 		  gnt_out_spec_qual;
		     assign gnt_out_spec_qual = |gnt_out_spec_qual_ip;
		     
		     assign sel_ip = gnt_out_nonspec_ip | gnt_out_spec_qual_ip;
		     
		     assign gnt = req_out_nonspec | gnt_out_spec_qual;
		     
		  end
		
	     end
	   else
	     begin
		assign gnt_out_spec_ip = {num_ports{1'b0}};
		assign gnt = req_out_nonspec;
		assign sel_ip = gnt_out_nonspec_ip;
	     end
	   
	   wire [0:num_vcs-1] sel_ivc;
	   c_select_1ofn
	     #(.num_ports(num_ports),
	       .width(num_vcs))
	   sel_ivc_sel
	     (.select(sel_ip),
	      .data_in(sel_ip_ivc),
	      .data_out(sel_ivc));
	   
	   assign gnt_out_nonspec_op_ip[op*num_ports:(op+1)*num_ports-1]
	     = gnt_out_nonspec_ip;
	   assign gnt_out_spec_op_ip[op*num_ports:(op+1)*num_ports-1]
	     = gnt_out_spec_ip;
	   assign gnt_op[op] = gnt;
	   assign sel_op_ip[op*num_ports:(op+1)*num_ports-1] = sel_ip;
	   assign sel_op_ivc[op*num_vcs:(op+1)*num_vcs-1] = sel_ivc;
	   
	end
      
   endgenerate
   
endmodule
