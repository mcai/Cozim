// $Id: c_fbgen.v 5188 2012-08-30 00:31:31Z dub $

/*
 Copyright (c) 2007-2012, Trustees of The Leland Stanford Junior University
 All rights reserved.

 Redistribution and use in source and binary forms, with or without
 modification, are permitted provided that the following conditions are met:

 Redistributions of source code must retain the above copyright notice, this 
 list of conditions and the following disclaimer.
 Redistributions in binary form must reproduce the above copyright notice, this
 list of conditions and the following disclaimer in the documentation and/or
 other materials provided with the distribution.

 THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
 ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
 WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE 
 DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR
 ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
 (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
 LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON
 ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
 (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
 SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/

//==============================================================================
// generic feedback polynomial generator
//==============================================================================

// NOTE: This file was automatically generated. Do not edit by hand!

module c_fbgen
  (feedback);
   
`include "c_constants.sv"
   
   // width of register (must be greater than one)
   parameter width = 32;
   
   // select one of possibly multiple provided polynomials
   parameter index = 0;
   
   // generated feedback polynomial
   output [0:width-1] feedback;
   wire [0:width-1] feedback;
   
   generate
      
      if(width == 1)
	begin
	   assign feedback = 1'h1;
	end
      else if(width == 2)
	begin
	   assign feedback = 2'h3;
	end
      else if(width == 3)
	begin
	   if((index % 2) == 0) assign feedback = 3'h5;
	   else if((index % 2) == 1) assign feedback = 3'h6;
	end
      else if(width == 4)
         begin
            if((index % 2) == 0) assign feedback = 4'h9;
            else if((index % 2) == 1) assign feedback = 4'hC;
         end
      else if(width == 5)
         begin
            if((index % 6) == 0) assign feedback = 5'h12;
            else if((index % 6) == 1) assign feedback = 5'h14;
            else if((index % 6) == 2) assign feedback = 5'h17;
            else if((index % 6) == 3) assign feedback = 5'h1B;
            else if((index % 6) == 4) assign feedback = 5'h1D;
            else if((index % 6) == 5) assign feedback = 5'h1E;
         end
      else if(width == 6)
         begin
            if((index % 6) == 0) assign feedback = 6'h21;
            else if((index % 6) == 1) assign feedback = 6'h2D;
            else if((index % 6) == 2) assign feedback = 6'h30;
            else if((index % 6) == 3) assign feedback = 6'h33;
            else if((index % 6) == 4) assign feedback = 6'h36;
            else if((index % 6) == 5) assign feedback = 6'h39;
         end
      else if(width == 7)
         begin
            if((index % 18) == 0) assign feedback = 7'h41;
            else if((index % 18) == 1) assign feedback = 7'h44;
            else if((index % 18) == 2) assign feedback = 7'h47;
            else if((index % 18) == 3) assign feedback = 7'h48;
            else if((index % 18) == 4) assign feedback = 7'h4E;
            else if((index % 18) == 5) assign feedback = 7'h53;
            else if((index % 18) == 6) assign feedback = 7'h55;
            else if((index % 18) == 7) assign feedback = 7'h5C;
            else if((index % 18) == 8) assign feedback = 7'h5F;
            else if((index % 18) == 9) assign feedback = 7'h60;
            else if((index % 18) == 10) assign feedback = 7'h65;
            else if((index % 18) == 11) assign feedback = 7'h69;
            else if((index % 18) == 12) assign feedback = 7'h6A;
            else if((index % 18) == 13) assign feedback = 7'h72;
            else if((index % 18) == 14) assign feedback = 7'h77;
            else if((index % 18) == 15) assign feedback = 7'h78;
            else if((index % 18) == 16) assign feedback = 7'h7B;
            else if((index % 18) == 17) assign feedback = 7'h7E;
         end
      else if(width == 8)
         begin
            if((index % 16) == 0) assign feedback = 8'h8E;
            else if((index % 16) == 1) assign feedback = 8'h95;
            else if((index % 16) == 2) assign feedback = 8'h96;
            else if((index % 16) == 3) assign feedback = 8'hA6;
            else if((index % 16) == 4) assign feedback = 8'hAF;
            else if((index % 16) == 5) assign feedback = 8'hB1;
            else if((index % 16) == 6) assign feedback = 8'hB2;
            else if((index % 16) == 7) assign feedback = 8'hB4;
            else if((index % 16) == 8) assign feedback = 8'hB8;
            else if((index % 16) == 9) assign feedback = 8'hC3;
            else if((index % 16) == 10) assign feedback = 8'hC6;
            else if((index % 16) == 11) assign feedback = 8'hD4;
            else if((index % 16) == 12) assign feedback = 8'hE1;
            else if((index % 16) == 13) assign feedback = 8'hE7;
            else if((index % 16) == 14) assign feedback = 8'hF3;
            else if((index % 16) == 15) assign feedback = 8'hFA;
         end
      else if(width == 9)
         begin
            if((index % 48) == 0) assign feedback = 9'h108;
            else if((index % 48) == 1) assign feedback = 9'h10D;
            else if((index % 48) == 2) assign feedback = 9'h110;
            else if((index % 48) == 3) assign feedback = 9'h116;
            else if((index % 48) == 4) assign feedback = 9'h119;
            else if((index % 48) == 5) assign feedback = 9'h12C;
            else if((index % 48) == 6) assign feedback = 9'h12F;
            else if((index % 48) == 7) assign feedback = 9'h134;
            else if((index % 48) == 8) assign feedback = 9'h137;
            else if((index % 48) == 9) assign feedback = 9'h13B;
            else if((index % 48) == 10) assign feedback = 9'h13E;
            else if((index % 48) == 11) assign feedback = 9'h143;
            else if((index % 48) == 12) assign feedback = 9'h14A;
            else if((index % 48) == 13) assign feedback = 9'h151;
            else if((index % 48) == 14) assign feedback = 9'h152;
            else if((index % 48) == 15) assign feedback = 9'h157;
            else if((index % 48) == 16) assign feedback = 9'h15B;
            else if((index % 48) == 17) assign feedback = 9'h15E;
            else if((index % 48) == 18) assign feedback = 9'h167;
            else if((index % 48) == 19) assign feedback = 9'h168;
            else if((index % 48) == 20) assign feedback = 9'h16D;
            else if((index % 48) == 21) assign feedback = 9'h17A;
            else if((index % 48) == 22) assign feedback = 9'h17C;
            else if((index % 48) == 23) assign feedback = 9'h189;
            else if((index % 48) == 24) assign feedback = 9'h18A;
            else if((index % 48) == 25) assign feedback = 9'h18F;
            else if((index % 48) == 26) assign feedback = 9'h191;
            else if((index % 48) == 27) assign feedback = 9'h198;
            else if((index % 48) == 28) assign feedback = 9'h19D;
            else if((index % 48) == 29) assign feedback = 9'h1A7;
            else if((index % 48) == 30) assign feedback = 9'h1AD;
            else if((index % 48) == 31) assign feedback = 9'h1B0;
            else if((index % 48) == 32) assign feedback = 9'h1B5;
            else if((index % 48) == 33) assign feedback = 9'h1B6;
            else if((index % 48) == 34) assign feedback = 9'h1B9;
            else if((index % 48) == 35) assign feedback = 9'h1BF;
            else if((index % 48) == 36) assign feedback = 9'h1C2;
            else if((index % 48) == 37) assign feedback = 9'h1C7;
            else if((index % 48) == 38) assign feedback = 9'h1DA;
            else if((index % 48) == 39) assign feedback = 9'h1DC;
            else if((index % 48) == 40) assign feedback = 9'h1E3;
            else if((index % 48) == 41) assign feedback = 9'h1E5;
            else if((index % 48) == 42) assign feedback = 9'h1E6;
            else if((index % 48) == 43) assign feedback = 9'h1EA;
            else if((index % 48) == 44) assign feedback = 9'h1EC;
            else if((index % 48) == 45) assign feedback = 9'h1F1;
            else if((index % 48) == 46) assign feedback = 9'h1F4;
            else if((index % 48) == 47) assign feedback = 9'h1FD;
         end
      else if(width == 10)
         begin
            if((index % 60) == 0) assign feedback = 10'h204;
            else if((index % 60) == 1) assign feedback = 10'h20D;
            else if((index % 60) == 2) assign feedback = 10'h213;
            else if((index % 60) == 3) assign feedback = 10'h216;
            else if((index % 60) == 4) assign feedback = 10'h232;
            else if((index % 60) == 5) assign feedback = 10'h237;
            else if((index % 60) == 6) assign feedback = 10'h240;
            else if((index % 60) == 7) assign feedback = 10'h245;
            else if((index % 60) == 8) assign feedback = 10'h262;
            else if((index % 60) == 9) assign feedback = 10'h26B;
            else if((index % 60) == 10) assign feedback = 10'h273;
            else if((index % 60) == 11) assign feedback = 10'h279;
            else if((index % 60) == 12) assign feedback = 10'h27F;
            else if((index % 60) == 13) assign feedback = 10'h286;
            else if((index % 60) == 14) assign feedback = 10'h28C;
            else if((index % 60) == 15) assign feedback = 10'h291;
            else if((index % 60) == 16) assign feedback = 10'h298;
            else if((index % 60) == 17) assign feedback = 10'h29E;
            else if((index % 60) == 18) assign feedback = 10'h2A1;
            else if((index % 60) == 19) assign feedback = 10'h2AB;
            else if((index % 60) == 20) assign feedback = 10'h2B5;
            else if((index % 60) == 21) assign feedback = 10'h2C2;
            else if((index % 60) == 22) assign feedback = 10'h2C7;
            else if((index % 60) == 23) assign feedback = 10'h2CB;
            else if((index % 60) == 24) assign feedback = 10'h2D0;
            else if((index % 60) == 25) assign feedback = 10'h2E3;
            else if((index % 60) == 26) assign feedback = 10'h2F2;
            else if((index % 60) == 27) assign feedback = 10'h2FB;
            else if((index % 60) == 28) assign feedback = 10'h2FD;
            else if((index % 60) == 29) assign feedback = 10'h309;
            else if((index % 60) == 30) assign feedback = 10'h30A;
            else if((index % 60) == 31) assign feedback = 10'h312;
            else if((index % 60) == 32) assign feedback = 10'h31B;
            else if((index % 60) == 33) assign feedback = 10'h321;
            else if((index % 60) == 34) assign feedback = 10'h327;
            else if((index % 60) == 35) assign feedback = 10'h32D;
            else if((index % 60) == 36) assign feedback = 10'h33C;
            else if((index % 60) == 37) assign feedback = 10'h33F;
            else if((index % 60) == 38) assign feedback = 10'h344;
            else if((index % 60) == 39) assign feedback = 10'h35A;
            else if((index % 60) == 40) assign feedback = 10'h360;
            else if((index % 60) == 41) assign feedback = 10'h369;
            else if((index % 60) == 42) assign feedback = 10'h36F;
            else if((index % 60) == 43) assign feedback = 10'h37E;
            else if((index % 60) == 44) assign feedback = 10'h38B;
            else if((index % 60) == 45) assign feedback = 10'h38E;
            else if((index % 60) == 46) assign feedback = 10'h390;
            else if((index % 60) == 47) assign feedback = 10'h39C;
            else if((index % 60) == 48) assign feedback = 10'h3A3;
            else if((index % 60) == 49) assign feedback = 10'h3A6;
            else if((index % 60) == 50) assign feedback = 10'h3AA;
            else if((index % 60) == 51) assign feedback = 10'h3AC;
            else if((index % 60) == 52) assign feedback = 10'h3B1;
            else if((index % 60) == 53) assign feedback = 10'h3BE;
            else if((index % 60) == 54) assign feedback = 10'h3C6;
            else if((index % 60) == 55) assign feedback = 10'h3C9;
            else if((index % 60) == 56) assign feedback = 10'h3D8;
            else if((index % 60) == 57) assign feedback = 10'h3ED;
            else if((index % 60) == 58) assign feedback = 10'h3F9;
            else if((index % 60) == 59) assign feedback = 10'h3FC;
         end
      else if(width == 11)
         begin
            if((index % 100) == 0) assign feedback = 11'h402;
            else if((index % 100) == 1) assign feedback = 11'h40B;
            else if((index % 100) == 2) assign feedback = 11'h415;
            else if((index % 100) == 3) assign feedback = 11'h416;
            else if((index % 100) == 4) assign feedback = 11'h423;
            else if((index % 100) == 5) assign feedback = 11'h431;
            else if((index % 100) == 6) assign feedback = 11'h432;
            else if((index % 100) == 7) assign feedback = 11'h438;
            else if((index % 100) == 8) assign feedback = 11'h43D;
            else if((index % 100) == 9) assign feedback = 11'h446;
            else if((index % 100) == 10) assign feedback = 11'h44A;
            else if((index % 100) == 11) assign feedback = 11'h44F;
            else if((index % 100) == 12) assign feedback = 11'h454;
            else if((index % 100) == 13) assign feedback = 11'h458;
            else if((index % 100) == 14) assign feedback = 11'h467;
            else if((index % 100) == 15) assign feedback = 11'h468;
            else if((index % 100) == 16) assign feedback = 11'h470;
            else if((index % 100) == 17) assign feedback = 11'h473;
            else if((index % 100) == 18) assign feedback = 11'h475;
            else if((index % 100) == 19) assign feedback = 11'h47A;
            else if((index % 100) == 20) assign feedback = 11'h486;
            else if((index % 100) == 21) assign feedback = 11'h489;
            else if((index % 100) == 22) assign feedback = 11'h492;
            else if((index % 100) == 23) assign feedback = 11'h494;
            else if((index % 100) == 24) assign feedback = 11'h49D;
            else if((index % 100) == 25) assign feedback = 11'h49E;
            else if((index % 100) == 26) assign feedback = 11'h4A2;
            else if((index % 100) == 27) assign feedback = 11'h4A4;
            else if((index % 100) == 28) assign feedback = 11'h4A8;
            else if((index % 100) == 29) assign feedback = 11'h4AD;
            else if((index % 100) == 30) assign feedback = 11'h4B9;
            else if((index % 100) == 31) assign feedback = 11'h4BA;
            else if((index % 100) == 32) assign feedback = 11'h4BF;
            else if((index % 100) == 33) assign feedback = 11'h4C1;
            else if((index % 100) == 34) assign feedback = 11'h4C7;
            else if((index % 100) == 35) assign feedback = 11'h4D5;
            else if((index % 100) == 36) assign feedback = 11'h4D6;
            else if((index % 100) == 37) assign feedback = 11'h4DC;
            else if((index % 100) == 38) assign feedback = 11'h4E3;
            else if((index % 100) == 39) assign feedback = 11'h4EC;
            else if((index % 100) == 40) assign feedback = 11'h4F2;
            else if((index % 100) == 41) assign feedback = 11'h4FB;
            else if((index % 100) == 42) assign feedback = 11'h500;
            else if((index % 100) == 43) assign feedback = 11'h503;
            else if((index % 100) == 44) assign feedback = 11'h509;
            else if((index % 100) == 45) assign feedback = 11'h50A;
            else if((index % 100) == 46) assign feedback = 11'h514;
            else if((index % 100) == 47) assign feedback = 11'h524;
            else if((index % 100) == 48) assign feedback = 11'h530;
            else if((index % 100) == 49) assign feedback = 11'h536;
            else if((index % 100) == 50) assign feedback = 11'h53C;
            else if((index % 100) == 51) assign feedback = 11'h53F;
            else if((index % 100) == 52) assign feedback = 11'h542;
            else if((index % 100) == 53) assign feedback = 11'h548;
            else if((index % 100) == 54) assign feedback = 11'h54E;
            else if((index % 100) == 55) assign feedback = 11'h553;
            else if((index % 100) == 56) assign feedback = 11'h555;
            else if((index % 100) == 57) assign feedback = 11'h559;
            else if((index % 100) == 58) assign feedback = 11'h55A;
            else if((index % 100) == 59) assign feedback = 11'h56A;
            else if((index % 100) == 60) assign feedback = 11'h56F;
            else if((index % 100) == 61) assign feedback = 11'h574;
            else if((index % 100) == 62) assign feedback = 11'h577;
            else if((index % 100) == 63) assign feedback = 11'h578;
            else if((index % 100) == 64) assign feedback = 11'h57D;
            else if((index % 100) == 65) assign feedback = 11'h581;
            else if((index % 100) == 66) assign feedback = 11'h584;
            else if((index % 100) == 67) assign feedback = 11'h588;
            else if((index % 100) == 68) assign feedback = 11'h599;
            else if((index % 100) == 69) assign feedback = 11'h59F;
            else if((index % 100) == 70) assign feedback = 11'h5A0;
            else if((index % 100) == 71) assign feedback = 11'h5A5;
            else if((index % 100) == 72) assign feedback = 11'h5AC;
            else if((index % 100) == 73) assign feedback = 11'h5AF;
            else if((index % 100) == 74) assign feedback = 11'h5B2;
            else if((index % 100) == 75) assign feedback = 11'h5B7;
            else if((index % 100) == 76) assign feedback = 11'h5BE;
            else if((index % 100) == 77) assign feedback = 11'h5C3;
            else if((index % 100) == 78) assign feedback = 11'h5C5;
            else if((index % 100) == 79) assign feedback = 11'h5C9;
            else if((index % 100) == 80) assign feedback = 11'h5CA;
            else if((index % 100) == 81) assign feedback = 11'h5D7;
            else if((index % 100) == 82) assign feedback = 11'h5DB;
            else if((index % 100) == 83) assign feedback = 11'h5DE;
            else if((index % 100) == 84) assign feedback = 11'h5E4;
            else if((index % 100) == 85) assign feedback = 11'h5ED;
            else if((index % 100) == 86) assign feedback = 11'h5EE;
            else if((index % 100) == 87) assign feedback = 11'h5F3;
            else if((index % 100) == 88) assign feedback = 11'h5F6;
            else if((index % 100) == 89) assign feedback = 11'h605;
            else if((index % 100) == 90) assign feedback = 11'h606;
            else if((index % 100) == 91) assign feedback = 11'h60C;
            else if((index % 100) == 92) assign feedback = 11'h60F;
            else if((index % 100) == 93) assign feedback = 11'h62B;
            else if((index % 100) == 94) assign feedback = 11'h630;
            else if((index % 100) == 95) assign feedback = 11'h635;
            else if((index % 100) == 96) assign feedback = 11'h639;
            else if((index % 100) == 97) assign feedback = 11'h642;
            else if((index % 100) == 98) assign feedback = 11'h644;
            else if((index % 100) == 99) assign feedback = 11'h64B;
         end
      else if(width == 12)
         begin
            if((index % 100) == 0) assign feedback = 12'h829;
            else if((index % 100) == 1) assign feedback = 12'h834;
            else if((index % 100) == 2) assign feedback = 12'h83D;
            else if((index % 100) == 3) assign feedback = 12'h83E;
            else if((index % 100) == 4) assign feedback = 12'h84C;
            else if((index % 100) == 5) assign feedback = 12'h868;
            else if((index % 100) == 6) assign feedback = 12'h875;
            else if((index % 100) == 7) assign feedback = 12'h883;
            else if((index % 100) == 8) assign feedback = 12'h88F;
            else if((index % 100) == 9) assign feedback = 12'h891;
            else if((index % 100) == 10) assign feedback = 12'h89D;
            else if((index % 100) == 11) assign feedback = 12'h8A7;
            else if((index % 100) == 12) assign feedback = 12'h8AB;
            else if((index % 100) == 13) assign feedback = 12'h8B0;
            else if((index % 100) == 14) assign feedback = 12'h8B5;
            else if((index % 100) == 15) assign feedback = 12'h8C2;
            else if((index % 100) == 16) assign feedback = 12'h8D9;
            else if((index % 100) == 17) assign feedback = 12'h8EC;
            else if((index % 100) == 18) assign feedback = 12'h8EF;
            else if((index % 100) == 19) assign feedback = 12'h906;
            else if((index % 100) == 20) assign feedback = 12'h91B;
            else if((index % 100) == 21) assign feedback = 12'h91E;
            else if((index % 100) == 22) assign feedback = 12'h933;
            else if((index % 100) == 23) assign feedback = 12'h939;
            else if((index % 100) == 24) assign feedback = 12'h93F;
            else if((index % 100) == 25) assign feedback = 12'h95C;
            else if((index % 100) == 26) assign feedback = 12'h960;
            else if((index % 100) == 27) assign feedback = 12'h965;
            else if((index % 100) == 28) assign feedback = 12'h987;
            else if((index % 100) == 29) assign feedback = 12'h98E;
            else if((index % 100) == 30) assign feedback = 12'h990;
            else if((index % 100) == 31) assign feedback = 12'h99C;
            else if((index % 100) == 32) assign feedback = 12'h99F;
            else if((index % 100) == 33) assign feedback = 12'h9A6;
            else if((index % 100) == 34) assign feedback = 12'h9B8;
            else if((index % 100) == 35) assign feedback = 12'h9CC;
            else if((index % 100) == 36) assign feedback = 12'h9D1;
            else if((index % 100) == 37) assign feedback = 12'h9D4;
            else if((index % 100) == 38) assign feedback = 12'hA03;
            else if((index % 100) == 39) assign feedback = 12'hA18;
            else if((index % 100) == 40) assign feedback = 12'hA1B;
            else if((index % 100) == 41) assign feedback = 12'hA27;
            else if((index % 100) == 42) assign feedback = 12'hA2E;
            else if((index % 100) == 43) assign feedback = 12'hA33;
            else if((index % 100) == 44) assign feedback = 12'hA3A;
            else if((index % 100) == 45) assign feedback = 12'hA53;
            else if((index % 100) == 46) assign feedback = 12'hA56;
            else if((index % 100) == 47) assign feedback = 12'hA69;
            else if((index % 100) == 48) assign feedback = 12'hA87;
            else if((index % 100) == 49) assign feedback = 12'hA8E;
            else if((index % 100) == 50) assign feedback = 12'hAA6;
            else if((index % 100) == 51) assign feedback = 12'hAC9;
            else if((index % 100) == 52) assign feedback = 12'hAE2;
            else if((index % 100) == 53) assign feedback = 12'hAEB;
            else if((index % 100) == 54) assign feedback = 12'hAEE;
            else if((index % 100) == 55) assign feedback = 12'hAF5;
            else if((index % 100) == 56) assign feedback = 12'hB04;
            else if((index % 100) == 57) assign feedback = 12'hB23;
            else if((index % 100) == 58) assign feedback = 12'hB2A;
            else if((index % 100) == 59) assign feedback = 12'hB2C;
            else if((index % 100) == 60) assign feedback = 12'hB52;
            else if((index % 100) == 61) assign feedback = 12'hB5E;
            else if((index % 100) == 62) assign feedback = 12'hB8A;
            else if((index % 100) == 63) assign feedback = 12'hB8C;
            else if((index % 100) == 64) assign feedback = 12'hBA1;
            else if((index % 100) == 65) assign feedback = 12'hBA2;
            else if((index % 100) == 66) assign feedback = 12'hBBA;
            else if((index % 100) == 67) assign feedback = 12'hBC4;
            else if((index % 100) == 68) assign feedback = 12'hBD6;
            else if((index % 100) == 69) assign feedback = 12'hBD9;
            else if((index % 100) == 70) assign feedback = 12'hBDF;
            else if((index % 100) == 71) assign feedback = 12'hBE0;
            else if((index % 100) == 72) assign feedback = 12'hC2B;
            else if((index % 100) == 73) assign feedback = 12'hC2E;
            else if((index % 100) == 74) assign feedback = 12'hC48;
            else if((index % 100) == 75) assign feedback = 12'hC4B;
            else if((index % 100) == 76) assign feedback = 12'hC5C;
            else if((index % 100) == 77) assign feedback = 12'hC77;
            else if((index % 100) == 78) assign feedback = 12'hC8D;
            else if((index % 100) == 79) assign feedback = 12'hC9A;
            else if((index % 100) == 80) assign feedback = 12'hCA0;
            else if((index % 100) == 81) assign feedback = 12'hCB2;
            else if((index % 100) == 82) assign feedback = 12'hCBD;
            else if((index % 100) == 83) assign feedback = 12'hCC5;
            else if((index % 100) == 84) assign feedback = 12'hCD8;
            else if((index % 100) == 85) assign feedback = 12'hCDE;
            else if((index % 100) == 86) assign feedback = 12'hCE4;
            else if((index % 100) == 87) assign feedback = 12'hCE7;
            else if((index % 100) == 88) assign feedback = 12'hCF3;
            else if((index % 100) == 89) assign feedback = 12'hD0D;
            else if((index % 100) == 90) assign feedback = 12'hD15;
            else if((index % 100) == 91) assign feedback = 12'hD19;
            else if((index % 100) == 92) assign feedback = 12'hD34;
            else if((index % 100) == 93) assign feedback = 12'hD45;
            else if((index % 100) == 94) assign feedback = 12'hD68;
            else if((index % 100) == 95) assign feedback = 12'hD70;
            else if((index % 100) == 96) assign feedback = 12'hD7A;
            else if((index % 100) == 97) assign feedback = 12'hD85;
            else if((index % 100) == 98) assign feedback = 12'hD89;
            else if((index % 100) == 99) assign feedback = 12'hD8F;
         end
      else if(width == 13)
         begin
            if((index % 100) == 0) assign feedback = 13'h100D;
            else if((index % 100) == 1) assign feedback = 13'h1013;
            else if((index % 100) == 2) assign feedback = 13'h101A;
            else if((index % 100) == 3) assign feedback = 13'h1029;
            else if((index % 100) == 4) assign feedback = 13'h1032;
            else if((index % 100) == 5) assign feedback = 13'h1037;
            else if((index % 100) == 6) assign feedback = 13'h1045;
            else if((index % 100) == 7) assign feedback = 13'h1046;
            else if((index % 100) == 8) assign feedback = 13'h104F;
            else if((index % 100) == 9) assign feedback = 13'h1052;
            else if((index % 100) == 10) assign feedback = 13'h1057;
            else if((index % 100) == 11) assign feedback = 13'h105D;
            else if((index % 100) == 12) assign feedback = 13'h105E;
            else if((index % 100) == 13) assign feedback = 13'h1061;
            else if((index % 100) == 14) assign feedback = 13'h1064;
            else if((index % 100) == 15) assign feedback = 13'h1070;
            else if((index % 100) == 16) assign feedback = 13'h1079;
            else if((index % 100) == 17) assign feedback = 13'h1086;
            else if((index % 100) == 18) assign feedback = 13'h108A;
            else if((index % 100) == 19) assign feedback = 13'h1094;
            else if((index % 100) == 20) assign feedback = 13'h1097;
            else if((index % 100) == 21) assign feedback = 13'h109D;
            else if((index % 100) == 22) assign feedback = 13'h10A1;
            else if((index % 100) == 23) assign feedback = 13'h10B3;
            else if((index % 100) == 24) assign feedback = 13'h10B5;
            else if((index % 100) == 25) assign feedback = 13'h10BC;
            else if((index % 100) == 26) assign feedback = 13'h10C4;
            else if((index % 100) == 27) assign feedback = 13'h10CB;
            else if((index % 100) == 28) assign feedback = 13'h10CE;
            else if((index % 100) == 29) assign feedback = 13'h10DF;
            else if((index % 100) == 30) assign feedback = 13'h10E0;
            else if((index % 100) == 31) assign feedback = 13'h10E3;
            else if((index % 100) == 32) assign feedback = 13'h10E6;
            else if((index % 100) == 33) assign feedback = 13'h10EF;
            else if((index % 100) == 34) assign feedback = 13'h10F1;
            else if((index % 100) == 35) assign feedback = 13'h10F8;
            else if((index % 100) == 36) assign feedback = 13'h10FD;
            else if((index % 100) == 37) assign feedback = 13'h110C;
            else if((index % 100) == 38) assign feedback = 13'h1112;
            else if((index % 100) == 39) assign feedback = 13'h111B;
            else if((index % 100) == 40) assign feedback = 13'h111E;
            else if((index % 100) == 41) assign feedback = 13'h1121;
            else if((index % 100) == 42) assign feedback = 13'h112D;
            else if((index % 100) == 43) assign feedback = 13'h112E;
            else if((index % 100) == 44) assign feedback = 13'h113C;
            else if((index % 100) == 45) assign feedback = 13'h113F;
            else if((index % 100) == 46) assign feedback = 13'h1144;
            else if((index % 100) == 47) assign feedback = 13'h114B;
            else if((index % 100) == 48) assign feedback = 13'h114D;
            else if((index % 100) == 49) assign feedback = 13'h1159;
            else if((index % 100) == 50) assign feedback = 13'h115F;
            else if((index % 100) == 51) assign feedback = 13'h1166;
            else if((index % 100) == 52) assign feedback = 13'h1177;
            else if((index % 100) == 53) assign feedback = 13'h117B;
            else if((index % 100) == 54) assign feedback = 13'h117D;
            else if((index % 100) == 55) assign feedback = 13'h1182;
            else if((index % 100) == 56) assign feedback = 13'h1193;
            else if((index % 100) == 57) assign feedback = 13'h1195;
            else if((index % 100) == 58) assign feedback = 13'h11A3;
            else if((index % 100) == 59) assign feedback = 13'h11AA;
            else if((index % 100) == 60) assign feedback = 13'h11AC;
            else if((index % 100) == 61) assign feedback = 13'h11B7;
            else if((index % 100) == 62) assign feedback = 13'h11B8;
            else if((index % 100) == 63) assign feedback = 13'h11BE;
            else if((index % 100) == 64) assign feedback = 13'h11C3;
            else if((index % 100) == 65) assign feedback = 13'h11C6;
            else if((index % 100) == 66) assign feedback = 13'h11CA;
            else if((index % 100) == 67) assign feedback = 13'h11D1;
            else if((index % 100) == 68) assign feedback = 13'h11D4;
            else if((index % 100) == 69) assign feedback = 13'h11D8;
            else if((index % 100) == 70) assign feedback = 13'h11DB;
            else if((index % 100) == 71) assign feedback = 13'h11DD;
            else if((index % 100) == 72) assign feedback = 13'h11F0;
            else if((index % 100) == 73) assign feedback = 13'h11F6;
            else if((index % 100) == 74) assign feedback = 13'h11FC;
            else if((index % 100) == 75) assign feedback = 13'h1205;
            else if((index % 100) == 76) assign feedback = 13'h1209;
            else if((index % 100) == 77) assign feedback = 13'h120F;
            else if((index % 100) == 78) assign feedback = 13'h1212;
            else if((index % 100) == 79) assign feedback = 13'h1214;
            else if((index % 100) == 80) assign feedback = 13'h121E;
            else if((index % 100) == 81) assign feedback = 13'h1228;
            else if((index % 100) == 82) assign feedback = 13'h122B;
            else if((index % 100) == 83) assign feedback = 13'h1230;
            else if((index % 100) == 84) assign feedback = 13'h1236;
            else if((index % 100) == 85) assign feedback = 13'h123F;
            else if((index % 100) == 86) assign feedback = 13'h1241;
            else if((index % 100) == 87) assign feedback = 13'h124D;
            else if((index % 100) == 88) assign feedback = 13'h124E;
            else if((index % 100) == 89) assign feedback = 13'h125A;
            else if((index % 100) == 90) assign feedback = 13'h125F;
            else if((index % 100) == 91) assign feedback = 13'h1260;
            else if((index % 100) == 92) assign feedback = 13'h1263;
            else if((index % 100) == 93) assign feedback = 13'h1265;
            else if((index % 100) == 94) assign feedback = 13'h1271;
            else if((index % 100) == 95) assign feedback = 13'h1284;
            else if((index % 100) == 96) assign feedback = 13'h128B;
            else if((index % 100) == 97) assign feedback = 13'h128E;
            else if((index % 100) == 98) assign feedback = 13'h1290;
            else if((index % 100) == 99) assign feedback = 13'h1296;
         end
      else if(width == 14)
         begin
            if((index % 100) == 0) assign feedback = 14'h2015;
            else if((index % 100) == 1) assign feedback = 14'h201C;
            else if((index % 100) == 2) assign feedback = 14'h2029;
            else if((index % 100) == 3) assign feedback = 14'h202F;
            else if((index % 100) == 4) assign feedback = 14'h203D;
            else if((index % 100) == 5) assign feedback = 14'h2054;
            else if((index % 100) == 6) assign feedback = 14'h2057;
            else if((index % 100) == 7) assign feedback = 14'h205D;
            else if((index % 100) == 8) assign feedback = 14'h205E;
            else if((index % 100) == 9) assign feedback = 14'h2067;
            else if((index % 100) == 10) assign feedback = 14'h2075;
            else if((index % 100) == 11) assign feedback = 14'h2079;
            else if((index % 100) == 12) assign feedback = 14'h2086;
            else if((index % 100) == 13) assign feedback = 14'h2089;
            else if((index % 100) == 14) assign feedback = 14'h209D;
            else if((index % 100) == 15) assign feedback = 14'h20A1;
            else if((index % 100) == 16) assign feedback = 14'h20CD;
            else if((index % 100) == 17) assign feedback = 14'h20CE;
            else if((index % 100) == 18) assign feedback = 14'h20D3;
            else if((index % 100) == 19) assign feedback = 14'h20D6;
            else if((index % 100) == 20) assign feedback = 14'h20DA;
            else if((index % 100) == 21) assign feedback = 14'h20EA;
            else if((index % 100) == 22) assign feedback = 14'h20EC;
            else if((index % 100) == 23) assign feedback = 14'h20F8;
            else if((index % 100) == 24) assign feedback = 14'h2106;
            else if((index % 100) == 25) assign feedback = 14'h212B;
            else if((index % 100) == 26) assign feedback = 14'h2130;
            else if((index % 100) == 27) assign feedback = 14'h213F;
            else if((index % 100) == 28) assign feedback = 14'h2142;
            else if((index % 100) == 29) assign feedback = 14'h214E;
            else if((index % 100) == 30) assign feedback = 14'h2163;
            else if((index % 100) == 31) assign feedback = 14'h2165;
            else if((index % 100) == 32) assign feedback = 14'h2166;
            else if((index % 100) == 33) assign feedback = 14'h2171;
            else if((index % 100) == 34) assign feedback = 14'h2174;
            else if((index % 100) == 35) assign feedback = 14'h2177;
            else if((index % 100) == 36) assign feedback = 14'h2184;
            else if((index % 100) == 37) assign feedback = 14'h2190;
            else if((index % 100) == 38) assign feedback = 14'h219F;
            else if((index % 100) == 39) assign feedback = 14'h21BE;
            else if((index % 100) == 40) assign feedback = 14'h21C3;
            else if((index % 100) == 41) assign feedback = 14'h21CA;
            else if((index % 100) == 42) assign feedback = 14'h21D7;
            else if((index % 100) == 43) assign feedback = 14'h21E4;
            else if((index % 100) == 44) assign feedback = 14'h21F5;
            else if((index % 100) == 45) assign feedback = 14'h21F6;
            else if((index % 100) == 46) assign feedback = 14'h2205;
            else if((index % 100) == 47) assign feedback = 14'h2221;
            else if((index % 100) == 48) assign feedback = 14'h2239;
            else if((index % 100) == 49) assign feedback = 14'h2269;
            else if((index % 100) == 50) assign feedback = 14'h226A;
            else if((index % 100) == 51) assign feedback = 14'h226F;
            else if((index % 100) == 52) assign feedback = 14'h2271;
            else if((index % 100) == 53) assign feedback = 14'h227D;
            else if((index % 100) == 54) assign feedback = 14'h2295;
            else if((index % 100) == 55) assign feedback = 14'h229C;
            else if((index % 100) == 56) assign feedback = 14'h22AC;
            else if((index % 100) == 57) assign feedback = 14'h22B7;
            else if((index % 100) == 58) assign feedback = 14'h22CC;
            else if((index % 100) == 59) assign feedback = 14'h22CF;
            else if((index % 100) == 60) assign feedback = 14'h22D2;
            else if((index % 100) == 61) assign feedback = 14'h22DB;
            else if((index % 100) == 62) assign feedback = 14'h22E2;
            else if((index % 100) == 63) assign feedback = 14'h22EB;
            else if((index % 100) == 64) assign feedback = 14'h22F3;
            else if((index % 100) == 65) assign feedback = 14'h22F9;
            else if((index % 100) == 66) assign feedback = 14'h22FF;
            else if((index % 100) == 67) assign feedback = 14'h2307;
            else if((index % 100) == 68) assign feedback = 14'h230E;
            else if((index % 100) == 69) assign feedback = 14'h2313;
            else if((index % 100) == 70) assign feedback = 14'h231A;
            else if((index % 100) == 71) assign feedback = 14'h2323;
            else if((index % 100) == 72) assign feedback = 14'h232C;
            else if((index % 100) == 73) assign feedback = 14'h2331;
            else if((index % 100) == 74) assign feedback = 14'h2338;
            else if((index % 100) == 75) assign feedback = 14'h233D;
            else if((index % 100) == 76) assign feedback = 14'h2352;
            else if((index % 100) == 77) assign feedback = 14'h2362;
            else if((index % 100) == 78) assign feedback = 14'h2367;
            else if((index % 100) == 79) assign feedback = 14'h236D;
            else if((index % 100) == 80) assign feedback = 14'h2398;
            else if((index % 100) == 81) assign feedback = 14'h23A7;
            else if((index % 100) == 82) assign feedback = 14'h23BF;
            else if((index % 100) == 83) assign feedback = 14'h23D3;
            else if((index % 100) == 84) assign feedback = 14'h23E0;
            else if((index % 100) == 85) assign feedback = 14'h23F2;
            else if((index % 100) == 86) assign feedback = 14'h23F4;
            else if((index % 100) == 87) assign feedback = 14'h23F7;
            else if((index % 100) == 88) assign feedback = 14'h2409;
            else if((index % 100) == 89) assign feedback = 14'h240C;
            else if((index % 100) == 90) assign feedback = 14'h241D;
            else if((index % 100) == 91) assign feedback = 14'h2421;
            else if((index % 100) == 92) assign feedback = 14'h242D;
            else if((index % 100) == 93) assign feedback = 14'h2430;
            else if((index % 100) == 94) assign feedback = 14'h2433;
            else if((index % 100) == 95) assign feedback = 14'h243F;
            else if((index % 100) == 96) assign feedback = 14'h2441;
            else if((index % 100) == 97) assign feedback = 14'h2471;
            else if((index % 100) == 98) assign feedback = 14'h248E;
            else if((index % 100) == 99) assign feedback = 14'h2496;
         end
      else if(width == 15)
         begin
            if((index % 100) == 0) assign feedback = 15'h4001;
            else if((index % 100) == 1) assign feedback = 15'h4008;
            else if((index % 100) == 2) assign feedback = 15'h400B;
            else if((index % 100) == 3) assign feedback = 15'h4016;
            else if((index % 100) == 4) assign feedback = 15'h401A;
            else if((index % 100) == 5) assign feedback = 15'h402F;
            else if((index % 100) == 6) assign feedback = 15'h403B;
            else if((index % 100) == 7) assign feedback = 15'h4040;
            else if((index % 100) == 8) assign feedback = 15'h4043;
            else if((index % 100) == 9) assign feedback = 15'h4049;
            else if((index % 100) == 10) assign feedback = 15'h4052;
            else if((index % 100) == 11) assign feedback = 15'h4061;
            else if((index % 100) == 12) assign feedback = 15'h4067;
            else if((index % 100) == 13) assign feedback = 15'h406E;
            else if((index % 100) == 14) assign feedback = 15'h4073;
            else if((index % 100) == 15) assign feedback = 15'h407A;
            else if((index % 100) == 16) assign feedback = 15'h4080;
            else if((index % 100) == 17) assign feedback = 15'h408A;
            else if((index % 100) == 18) assign feedback = 15'h4092;
            else if((index % 100) == 19) assign feedback = 15'h40AB;
            else if((index % 100) == 20) assign feedback = 15'h40AE;
            else if((index % 100) == 21) assign feedback = 15'h40B0;
            else if((index % 100) == 22) assign feedback = 15'h40B6;
            else if((index % 100) == 23) assign feedback = 15'h40C2;
            else if((index % 100) == 24) assign feedback = 15'h40D0;
            else if((index % 100) == 25) assign feedback = 15'h40D3;
            else if((index % 100) == 26) assign feedback = 15'h40DC;
            else if((index % 100) == 27) assign feedback = 15'h40E5;
            else if((index % 100) == 28) assign feedback = 15'h40E6;
            else if((index % 100) == 29) assign feedback = 15'h40EF;
            else if((index % 100) == 30) assign feedback = 15'h40FE;
            else if((index % 100) == 31) assign feedback = 15'h4109;
            else if((index % 100) == 32) assign feedback = 15'h411D;
            else if((index % 100) == 33) assign feedback = 15'h4122;
            else if((index % 100) == 34) assign feedback = 15'h413F;
            else if((index % 100) == 35) assign feedback = 15'h4144;
            else if((index % 100) == 36) assign feedback = 15'h4147;
            else if((index % 100) == 37) assign feedback = 15'h414D;
            else if((index % 100) == 38) assign feedback = 15'h4165;
            else if((index % 100) == 39) assign feedback = 15'h416C;
            else if((index % 100) == 40) assign feedback = 15'h418B;
            else if((index % 100) == 41) assign feedback = 15'h418D;
            else if((index % 100) == 42) assign feedback = 15'h4195;
            else if((index % 100) == 43) assign feedback = 15'h4199;
            else if((index % 100) == 44) assign feedback = 15'h41A3;
            else if((index % 100) == 45) assign feedback = 15'h41A6;
            else if((index % 100) == 46) assign feedback = 15'h41AF;
            else if((index % 100) == 47) assign feedback = 15'h41B1;
            else if((index % 100) == 48) assign feedback = 15'h41B4;
            else if((index % 100) == 49) assign feedback = 15'h41B8;
            else if((index % 100) == 50) assign feedback = 15'h41C5;
            else if((index % 100) == 51) assign feedback = 15'h41CC;
            else if((index % 100) == 52) assign feedback = 15'h41D7;
            else if((index % 100) == 53) assign feedback = 15'h41DE;
            else if((index % 100) == 54) assign feedback = 15'h41E2;
            else if((index % 100) == 55) assign feedback = 15'h41E8;
            else if((index % 100) == 56) assign feedback = 15'h420C;
            else if((index % 100) == 57) assign feedback = 15'h4211;
            else if((index % 100) == 58) assign feedback = 15'h4217;
            else if((index % 100) == 59) assign feedback = 15'h4218;
            else if((index % 100) == 60) assign feedback = 15'h421B;
            else if((index % 100) == 61) assign feedback = 15'h4233;
            else if((index % 100) == 62) assign feedback = 15'h4236;
            else if((index % 100) == 63) assign feedback = 15'h423C;
            else if((index % 100) == 64) assign feedback = 15'h4241;
            else if((index % 100) == 65) assign feedback = 15'h424B;
            else if((index % 100) == 66) assign feedback = 15'h4250;
            else if((index % 100) == 67) assign feedback = 15'h425A;
            else if((index % 100) == 68) assign feedback = 15'h426F;
            else if((index % 100) == 69) assign feedback = 15'h427B;
            else if((index % 100) == 70) assign feedback = 15'h427E;
            else if((index % 100) == 71) assign feedback = 15'h428E;
            else if((index % 100) == 72) assign feedback = 15'h4290;
            else if((index % 100) == 73) assign feedback = 15'h4293;
            else if((index % 100) == 74) assign feedback = 15'h4299;
            else if((index % 100) == 75) assign feedback = 15'h42A3;
            else if((index % 100) == 76) assign feedback = 15'h42A5;
            else if((index % 100) == 77) assign feedback = 15'h42AF;
            else if((index % 100) == 78) assign feedback = 15'h42B8;
            else if((index % 100) == 79) assign feedback = 15'h42BD;
            else if((index % 100) == 80) assign feedback = 15'h42C0;
            else if((index % 100) == 81) assign feedback = 15'h42C6;
            else if((index % 100) == 82) assign feedback = 15'h42D1;
            else if((index % 100) == 83) assign feedback = 15'h42D8;
            else if((index % 100) == 84) assign feedback = 15'h42E2;
            else if((index % 100) == 85) assign feedback = 15'h42E4;
            else if((index % 100) == 86) assign feedback = 15'h42ED;
            else if((index % 100) == 87) assign feedback = 15'h42F6;
            else if((index % 100) == 88) assign feedback = 15'h42F9;
            else if((index % 100) == 89) assign feedback = 15'h4304;
            else if((index % 100) == 90) assign feedback = 15'h4308;
            else if((index % 100) == 91) assign feedback = 15'h430E;
            else if((index % 100) == 92) assign feedback = 15'h4315;
            else if((index % 100) == 93) assign feedback = 15'h432A;
            else if((index % 100) == 94) assign feedback = 15'h432C;
            else if((index % 100) == 95) assign feedback = 15'h4332;
            else if((index % 100) == 96) assign feedback = 15'h433E;
            else if((index % 100) == 97) assign feedback = 15'h4340;
            else if((index % 100) == 98) assign feedback = 15'h4354;
            else if((index % 100) == 99) assign feedback = 15'h4357;
         end
      else if(width == 16)
         begin
            if((index % 100) == 0) assign feedback = 16'h8016;
            else if((index % 100) == 1) assign feedback = 16'h801C;
            else if((index % 100) == 2) assign feedback = 16'h801F;
            else if((index % 100) == 3) assign feedback = 16'h8029;
            else if((index % 100) == 4) assign feedback = 16'h805E;
            else if((index % 100) == 5) assign feedback = 16'h806B;
            else if((index % 100) == 6) assign feedback = 16'h8097;
            else if((index % 100) == 7) assign feedback = 16'h809E;
            else if((index % 100) == 8) assign feedback = 16'h80A7;
            else if((index % 100) == 9) assign feedback = 16'h80AE;
            else if((index % 100) == 10) assign feedback = 16'h80CB;
            else if((index % 100) == 11) assign feedback = 16'h80D0;
            else if((index % 100) == 12) assign feedback = 16'h80D6;
            else if((index % 100) == 13) assign feedback = 16'h80DF;
            else if((index % 100) == 14) assign feedback = 16'h80E3;
            else if((index % 100) == 15) assign feedback = 16'h810A;
            else if((index % 100) == 16) assign feedback = 16'h810C;
            else if((index % 100) == 17) assign feedback = 16'h8112;
            else if((index % 100) == 18) assign feedback = 16'h8117;
            else if((index % 100) == 19) assign feedback = 16'h812E;
            else if((index % 100) == 20) assign feedback = 16'h8136;
            else if((index % 100) == 21) assign feedback = 16'h8142;
            else if((index % 100) == 22) assign feedback = 16'h8148;
            else if((index % 100) == 23) assign feedback = 16'h8150;
            else if((index % 100) == 24) assign feedback = 16'h8172;
            else if((index % 100) == 25) assign feedback = 16'h818E;
            else if((index % 100) == 26) assign feedback = 16'h81A5;
            else if((index % 100) == 27) assign feedback = 16'h81B4;
            else if((index % 100) == 28) assign feedback = 16'h81B8;
            else if((index % 100) == 29) assign feedback = 16'h81C3;
            else if((index % 100) == 30) assign feedback = 16'h81C6;
            else if((index % 100) == 31) assign feedback = 16'h81CF;
            else if((index % 100) == 32) assign feedback = 16'h81D1;
            else if((index % 100) == 33) assign feedback = 16'h81EE;
            else if((index % 100) == 34) assign feedback = 16'h81FC;
            else if((index % 100) == 35) assign feedback = 16'h8214;
            else if((index % 100) == 36) assign feedback = 16'h822B;
            else if((index % 100) == 37) assign feedback = 16'h8233;
            else if((index % 100) == 38) assign feedback = 16'h8241;
            else if((index % 100) == 39) assign feedback = 16'h8244;
            else if((index % 100) == 40) assign feedback = 16'h8248;
            else if((index % 100) == 41) assign feedback = 16'h825F;
            else if((index % 100) == 42) assign feedback = 16'h8260;
            else if((index % 100) == 43) assign feedback = 16'h8299;
            else if((index % 100) == 44) assign feedback = 16'h82A3;
            else if((index % 100) == 45) assign feedback = 16'h82B4;
            else if((index % 100) == 46) assign feedback = 16'h82C3;
            else if((index % 100) == 47) assign feedback = 16'h82E1;
            else if((index % 100) == 48) assign feedback = 16'h82EE;
            else if((index % 100) == 49) assign feedback = 16'h82F5;
            else if((index % 100) == 50) assign feedback = 16'h8320;
            else if((index % 100) == 51) assign feedback = 16'h8325;
            else if((index % 100) == 52) assign feedback = 16'h8329;
            else if((index % 100) == 53) assign feedback = 16'h8345;
            else if((index % 100) == 54) assign feedback = 16'h8361;
            else if((index % 100) == 55) assign feedback = 16'h83B5;
            else if((index % 100) == 56) assign feedback = 16'h83B6;
            else if((index % 100) == 57) assign feedback = 16'h83BC;
            else if((index % 100) == 58) assign feedback = 16'h83C1;
            else if((index % 100) == 59) assign feedback = 16'h83F8;
            else if((index % 100) == 60) assign feedback = 16'h8406;
            else if((index % 100) == 61) assign feedback = 16'h8430;
            else if((index % 100) == 62) assign feedback = 16'h845F;
            else if((index % 100) == 63) assign feedback = 16'h846A;
            else if((index % 100) == 64) assign feedback = 16'h846F;
            else if((index % 100) == 65) assign feedback = 16'h8471;
            else if((index % 100) == 66) assign feedback = 16'h8478;
            else if((index % 100) == 67) assign feedback = 16'h847D;
            else if((index % 100) == 68) assign feedback = 16'h849C;
            else if((index % 100) == 69) assign feedback = 16'h84BE;
            else if((index % 100) == 70) assign feedback = 16'h84C5;
            else if((index % 100) == 71) assign feedback = 16'h84D2;
            else if((index % 100) == 72) assign feedback = 16'h84D7;
            else if((index % 100) == 73) assign feedback = 16'h84E1;
            else if((index % 100) == 74) assign feedback = 16'h84E2;
            else if((index % 100) == 75) assign feedback = 16'h84F3;
            else if((index % 100) == 76) assign feedback = 16'h84F9;
            else if((index % 100) == 77) assign feedback = 16'h853E;
            else if((index % 100) == 78) assign feedback = 16'h8540;
            else if((index % 100) == 79) assign feedback = 16'h855D;
            else if((index % 100) == 80) assign feedback = 16'h8562;
            else if((index % 100) == 81) assign feedback = 16'h8580;
            else if((index % 100) == 82) assign feedback = 16'h8589;
            else if((index % 100) == 83) assign feedback = 16'h858A;
            else if((index % 100) == 84) assign feedback = 16'h85A8;
            else if((index % 100) == 85) assign feedback = 16'h85AE;
            else if((index % 100) == 86) assign feedback = 16'h85E6;
            else if((index % 100) == 87) assign feedback = 16'h85E9;
            else if((index % 100) == 88) assign feedback = 16'h85F2;
            else if((index % 100) == 89) assign feedback = 16'h8607;
            else if((index % 100) == 90) assign feedback = 16'h860E;
            else if((index % 100) == 91) assign feedback = 16'h8610;
            else if((index % 100) == 92) assign feedback = 16'h8634;
            else if((index % 100) == 93) assign feedback = 16'h8638;
            else if((index % 100) == 94) assign feedback = 16'h863D;
            else if((index % 100) == 95) assign feedback = 16'h8646;
            else if((index % 100) == 96) assign feedback = 16'h864A;
            else if((index % 100) == 97) assign feedback = 16'h8651;
            else if((index % 100) == 98) assign feedback = 16'h8657;
            else if((index % 100) == 99) assign feedback = 16'h8679;
         end
      else if(width == 17)
         begin
            if((index % 100) == 0) assign feedback = 17'h10004;
            else if((index % 100) == 1) assign feedback = 17'h10007;
            else if((index % 100) == 2) assign feedback = 17'h10010;
            else if((index % 100) == 3) assign feedback = 17'h10016;
            else if((index % 100) == 4) assign feedback = 17'h10019;
            else if((index % 100) == 5) assign feedback = 17'h1001F;
            else if((index % 100) == 6) assign feedback = 17'h10020;
            else if((index % 100) == 7) assign feedback = 17'h1002A;
            else if((index % 100) == 8) assign feedback = 17'h10034;
            else if((index % 100) == 9) assign feedback = 17'h1003D;
            else if((index % 100) == 10) assign feedback = 17'h10046;
            else if((index % 100) == 11) assign feedback = 17'h1004C;
            else if((index % 100) == 12) assign feedback = 17'h10051;
            else if((index % 100) == 13) assign feedback = 17'h10057;
            else if((index % 100) == 14) assign feedback = 17'h1005D;
            else if((index % 100) == 15) assign feedback = 17'h10062;
            else if((index % 100) == 16) assign feedback = 17'h1007A;
            else if((index % 100) == 17) assign feedback = 17'h10085;
            else if((index % 100) == 18) assign feedback = 17'h10086;
            else if((index % 100) == 19) assign feedback = 17'h1008C;
            else if((index % 100) == 20) assign feedback = 17'h10092;
            else if((index % 100) == 21) assign feedback = 17'h1009E;
            else if((index % 100) == 22) assign feedback = 17'h100AB;
            else if((index % 100) == 23) assign feedback = 17'h100B0;
            else if((index % 100) == 24) assign feedback = 17'h100B3;
            else if((index % 100) == 25) assign feedback = 17'h100B6;
            else if((index % 100) == 26) assign feedback = 17'h100BF;
            else if((index % 100) == 27) assign feedback = 17'h100C1;
            else if((index % 100) == 28) assign feedback = 17'h100E0;
            else if((index % 100) == 29) assign feedback = 17'h100E3;
            else if((index % 100) == 30) assign feedback = 17'h100E5;
            else if((index % 100) == 31) assign feedback = 17'h100EC;
            else if((index % 100) == 32) assign feedback = 17'h100F8;
            else if((index % 100) == 33) assign feedback = 17'h10106;
            else if((index % 100) == 34) assign feedback = 17'h10111;
            else if((index % 100) == 35) assign feedback = 17'h10114;
            else if((index % 100) == 36) assign feedback = 17'h10118;
            else if((index % 100) == 37) assign feedback = 17'h1011B;
            else if((index % 100) == 38) assign feedback = 17'h10122;
            else if((index % 100) == 39) assign feedback = 17'h10135;
            else if((index % 100) == 40) assign feedback = 17'h1013C;
            else if((index % 100) == 41) assign feedback = 17'h1013F;
            else if((index % 100) == 42) assign feedback = 17'h10141;
            else if((index % 100) == 43) assign feedback = 17'h10148;
            else if((index % 100) == 44) assign feedback = 17'h1015A;
            else if((index % 100) == 45) assign feedback = 17'h10163;
            else if((index % 100) == 46) assign feedback = 17'h1016F;
            else if((index % 100) == 47) assign feedback = 17'h10171;
            else if((index % 100) == 48) assign feedback = 17'h10174;
            else if((index % 100) == 49) assign feedback = 17'h1017E;
            else if((index % 100) == 50) assign feedback = 17'h10184;
            else if((index % 100) == 51) assign feedback = 17'h10188;
            else if((index % 100) == 52) assign feedback = 17'h1018B;
            else if((index % 100) == 53) assign feedback = 17'h1018D;
            else if((index % 100) == 54) assign feedback = 17'h10193;
            else if((index % 100) == 55) assign feedback = 17'h10199;
            else if((index % 100) == 56) assign feedback = 17'h1019A;
            else if((index % 100) == 57) assign feedback = 17'h101A9;
            else if((index % 100) == 58) assign feedback = 17'h101BB;
            else if((index % 100) == 59) assign feedback = 17'h101D8;
            else if((index % 100) == 60) assign feedback = 17'h101DB;
            else if((index % 100) == 61) assign feedback = 17'h101E1;
            else if((index % 100) == 62) assign feedback = 17'h101E8;
            else if((index % 100) == 63) assign feedback = 17'h101ED;
            else if((index % 100) == 64) assign feedback = 17'h101F5;
            else if((index % 100) == 65) assign feedback = 17'h10203;
            else if((index % 100) == 66) assign feedback = 17'h1020A;
            else if((index % 100) == 67) assign feedback = 17'h1020C;
            else if((index % 100) == 68) assign feedback = 17'h1020F;
            else if((index % 100) == 69) assign feedback = 17'h10217;
            else if((index % 100) == 70) assign feedback = 17'h1021E;
            else if((index % 100) == 71) assign feedback = 17'h10221;
            else if((index % 100) == 72) assign feedback = 17'h1022B;
            else if((index % 100) == 73) assign feedback = 17'h1022E;
            else if((index % 100) == 74) assign feedback = 17'h10230;
            else if((index % 100) == 75) assign feedback = 17'h10233;
            else if((index % 100) == 76) assign feedback = 17'h1023A;
            else if((index % 100) == 77) assign feedback = 17'h10242;
            else if((index % 100) == 78) assign feedback = 17'h10247;
            else if((index % 100) == 79) assign feedback = 17'h1024E;
            else if((index % 100) == 80) assign feedback = 17'h10255;
            else if((index % 100) == 81) assign feedback = 17'h1025C;
            else if((index % 100) == 82) assign feedback = 17'h10260;
            else if((index % 100) == 83) assign feedback = 17'h10266;
            else if((index % 100) == 84) assign feedback = 17'h1027B;
            else if((index % 100) == 85) assign feedback = 17'h1027D;
            else if((index % 100) == 86) assign feedback = 17'h1028D;
            else if((index % 100) == 87) assign feedback = 17'h1028E;
            else if((index % 100) == 88) assign feedback = 17'h10293;
            else if((index % 100) == 89) assign feedback = 17'h1029A;
            else if((index % 100) == 90) assign feedback = 17'h1029F;
            else if((index % 100) == 91) assign feedback = 17'h102B1;
            else if((index % 100) == 92) assign feedback = 17'h102B2;
            else if((index % 100) == 93) assign feedback = 17'h102B7;
            else if((index % 100) == 94) assign feedback = 17'h102C9;
            else if((index % 100) == 95) assign feedback = 17'h102D2;
            else if((index % 100) == 96) assign feedback = 17'h102DD;
            else if((index % 100) == 97) assign feedback = 17'h102F6;
            else if((index % 100) == 98) assign feedback = 17'h10302;
            else if((index % 100) == 99) assign feedback = 17'h1030E;
         end
      else if(width == 18)
         begin
            if((index % 100) == 0) assign feedback = 18'h20013;
            else if((index % 100) == 1) assign feedback = 18'h2001F;
            else if((index % 100) == 2) assign feedback = 18'h20026;
            else if((index % 100) == 3) assign feedback = 18'h2003D;
            else if((index % 100) == 4) assign feedback = 18'h20040;
            else if((index % 100) == 5) assign feedback = 18'h2006D;
            else if((index % 100) == 6) assign feedback = 18'h20073;
            else if((index % 100) == 7) assign feedback = 18'h20076;
            else if((index % 100) == 8) assign feedback = 18'h20083;
            else if((index % 100) == 9) assign feedback = 18'h200A7;
            else if((index % 100) == 10) assign feedback = 18'h200C8;
            else if((index % 100) == 11) assign feedback = 18'h200F1;
            else if((index % 100) == 12) assign feedback = 18'h200F4;
            else if((index % 100) == 13) assign feedback = 18'h200F7;
            else if((index % 100) == 14) assign feedback = 18'h20105;
            else if((index % 100) == 15) assign feedback = 18'h20109;
            else if((index % 100) == 16) assign feedback = 18'h20130;
            else if((index % 100) == 17) assign feedback = 18'h2013A;
            else if((index % 100) == 18) assign feedback = 18'h20155;
            else if((index % 100) == 19) assign feedback = 18'h20178;
            else if((index % 100) == 20) assign feedback = 18'h2018B;
            else if((index % 100) == 21) assign feedback = 18'h20195;
            else if((index % 100) == 22) assign feedback = 18'h20196;
            else if((index % 100) == 23) assign feedback = 18'h201BB;
            else if((index % 100) == 24) assign feedback = 18'h201C3;
            else if((index % 100) == 25) assign feedback = 18'h201CA;
            else if((index % 100) == 26) assign feedback = 18'h201CC;
            else if((index % 100) == 27) assign feedback = 18'h201D4;
            else if((index % 100) == 28) assign feedback = 18'h201D8;
            else if((index % 100) == 29) assign feedback = 18'h201E2;
            else if((index % 100) == 30) assign feedback = 18'h201EB;
            else if((index % 100) == 31) assign feedback = 18'h201F0;
            else if((index % 100) == 32) assign feedback = 18'h2020C;
            else if((index % 100) == 33) assign feedback = 18'h20218;
            else if((index % 100) == 34) assign feedback = 18'h2021E;
            else if((index % 100) == 35) assign feedback = 18'h2022D;
            else if((index % 100) == 36) assign feedback = 18'h2023C;
            else if((index % 100) == 37) assign feedback = 18'h20244;
            else if((index % 100) == 38) assign feedback = 18'h20250;
            else if((index % 100) == 39) assign feedback = 18'h20290;
            else if((index % 100) == 40) assign feedback = 18'h202C9;
            else if((index % 100) == 41) assign feedback = 18'h202CF;
            else if((index % 100) == 42) assign feedback = 18'h202E2;
            else if((index % 100) == 43) assign feedback = 18'h202ED;
            else if((index % 100) == 44) assign feedback = 18'h202F0;
            else if((index % 100) == 45) assign feedback = 18'h202FF;
            else if((index % 100) == 46) assign feedback = 18'h20304;
            else if((index % 100) == 47) assign feedback = 18'h2030E;
            else if((index % 100) == 48) assign feedback = 18'h20315;
            else if((index % 100) == 49) assign feedback = 18'h2033E;
            else if((index % 100) == 50) assign feedback = 18'h20346;
            else if((index % 100) == 51) assign feedback = 18'h20394;
            else if((index % 100) == 52) assign feedback = 18'h20398;
            else if((index % 100) == 53) assign feedback = 18'h203A8;
            else if((index % 100) == 54) assign feedback = 18'h203DF;
            else if((index % 100) == 55) assign feedback = 18'h203E6;
            else if((index % 100) == 56) assign feedback = 18'h203F8;
            else if((index % 100) == 57) assign feedback = 18'h20400;
            else if((index % 100) == 58) assign feedback = 18'h2041D;
            else if((index % 100) == 59) assign feedback = 18'h20439;
            else if((index % 100) == 60) assign feedback = 18'h20442;
            else if((index % 100) == 61) assign feedback = 18'h20465;
            else if((index % 100) == 62) assign feedback = 18'h2046F;
            else if((index % 100) == 63) assign feedback = 18'h20477;
            else if((index % 100) == 64) assign feedback = 18'h2047E;
            else if((index % 100) == 65) assign feedback = 18'h20482;
            else if((index % 100) == 66) assign feedback = 18'h20493;
            else if((index % 100) == 67) assign feedback = 18'h20496;
            else if((index % 100) == 68) assign feedback = 18'h204B2;
            else if((index % 100) == 69) assign feedback = 18'h204BD;
            else if((index % 100) == 70) assign feedback = 18'h204C9;
            else if((index % 100) == 71) assign feedback = 18'h204D1;
            else if((index % 100) == 72) assign feedback = 18'h204D2;
            else if((index % 100) == 73) assign feedback = 18'h204E4;
            else if((index % 100) == 74) assign feedback = 18'h204E7;
            else if((index % 100) == 75) assign feedback = 18'h2050E;
            else if((index % 100) == 76) assign feedback = 18'h20545;
            else if((index % 100) == 77) assign feedback = 18'h2054A;
            else if((index % 100) == 78) assign feedback = 18'h20562;
            else if((index % 100) == 79) assign feedback = 18'h20567;
            else if((index % 100) == 80) assign feedback = 18'h2056B;
            else if((index % 100) == 81) assign feedback = 18'h20570;
            else if((index % 100) == 82) assign feedback = 18'h2057A;
            else if((index % 100) == 83) assign feedback = 18'h2058C;
            else if((index % 100) == 84) assign feedback = 18'h20594;
            else if((index % 100) == 85) assign feedback = 18'h2059D;
            else if((index % 100) == 86) assign feedback = 18'h205A8;
            else if((index % 100) == 87) assign feedback = 18'h205B3;
            else if((index % 100) == 88) assign feedback = 18'h205C1;
            else if((index % 100) == 89) assign feedback = 18'h205E3;
            else if((index % 100) == 90) assign feedback = 18'h205EC;
            else if((index % 100) == 91) assign feedback = 18'h205F8;
            else if((index % 100) == 92) assign feedback = 18'h20625;
            else if((index % 100) == 93) assign feedback = 18'h20638;
            else if((index % 100) == 94) assign feedback = 18'h2063D;
            else if((index % 100) == 95) assign feedback = 18'h20676;
            else if((index % 100) == 96) assign feedback = 18'h2067F;
            else if((index % 100) == 97) assign feedback = 18'h206C2;
            else if((index % 100) == 98) assign feedback = 18'h206CB;
            else if((index % 100) == 99) assign feedback = 18'h206CD;
         end
      else if(width == 19)
         begin
            if((index % 100) == 0) assign feedback = 19'h40013;
            else if((index % 100) == 1) assign feedback = 19'h4001F;
            else if((index % 100) == 2) assign feedback = 19'h40023;
            else if((index % 100) == 3) assign feedback = 19'h40029;
            else if((index % 100) == 4) assign feedback = 19'h4002C;
            else if((index % 100) == 5) assign feedback = 19'h40031;
            else if((index % 100) == 6) assign feedback = 19'h40037;
            else if((index % 100) == 7) assign feedback = 19'h4003E;
            else if((index % 100) == 8) assign feedback = 19'h40049;
            else if((index % 100) == 9) assign feedback = 19'h40057;
            else if((index % 100) == 10) assign feedback = 19'h40070;
            else if((index % 100) == 11) assign feedback = 19'h400A1;
            else if((index % 100) == 12) assign feedback = 19'h400B0;
            else if((index % 100) == 13) assign feedback = 19'h400B5;
            else if((index % 100) == 14) assign feedback = 19'h400BA;
            else if((index % 100) == 15) assign feedback = 19'h400C2;
            else if((index % 100) == 16) assign feedback = 19'h400CE;
            else if((index % 100) == 17) assign feedback = 19'h400D0;
            else if((index % 100) == 18) assign feedback = 19'h400D6;
            else if((index % 100) == 19) assign feedback = 19'h400D9;
            else if((index % 100) == 20) assign feedback = 19'h400DF;
            else if((index % 100) == 21) assign feedback = 19'h400E3;
            else if((index % 100) == 22) assign feedback = 19'h400E6;
            else if((index % 100) == 23) assign feedback = 19'h400EF;
            else if((index % 100) == 24) assign feedback = 19'h40105;
            else if((index % 100) == 25) assign feedback = 19'h40109;
            else if((index % 100) == 26) assign feedback = 19'h4010C;
            else if((index % 100) == 27) assign feedback = 19'h40112;
            else if((index % 100) == 28) assign feedback = 19'h40118;
            else if((index % 100) == 29) assign feedback = 19'h40127;
            else if((index % 100) == 30) assign feedback = 19'h40128;
            else if((index % 100) == 31) assign feedback = 19'h40135;
            else if((index % 100) == 32) assign feedback = 19'h40136;
            else if((index % 100) == 33) assign feedback = 19'h40141;
            else if((index % 100) == 34) assign feedback = 19'h40142;
            else if((index % 100) == 35) assign feedback = 19'h4014B;
            else if((index % 100) == 36) assign feedback = 19'h40150;
            else if((index % 100) == 37) assign feedback = 19'h40190;
            else if((index % 100) == 38) assign feedback = 19'h401A3;
            else if((index % 100) == 39) assign feedback = 19'h401B4;
            else if((index % 100) == 40) assign feedback = 19'h401B7;
            else if((index % 100) == 41) assign feedback = 19'h401CF;
            else if((index % 100) == 42) assign feedback = 19'h401D2;
            else if((index % 100) == 43) assign feedback = 19'h401D4;
            else if((index % 100) == 44) assign feedback = 19'h401E4;
            else if((index % 100) == 45) assign feedback = 19'h401EB;
            else if((index % 100) == 46) assign feedback = 19'h401ED;
            else if((index % 100) == 47) assign feedback = 19'h401EE;
            else if((index % 100) == 48) assign feedback = 19'h401F9;
            else if((index % 100) == 49) assign feedback = 19'h4021B;
            else if((index % 100) == 50) assign feedback = 19'h40228;
            else if((index % 100) == 51) assign feedback = 19'h4023A;
            else if((index % 100) == 52) assign feedback = 19'h4023F;
            else if((index % 100) == 53) assign feedback = 19'h40244;
            else if((index % 100) == 54) assign feedback = 19'h40248;
            else if((index % 100) == 55) assign feedback = 19'h4025A;
            else if((index % 100) == 56) assign feedback = 19'h4025C;
            else if((index % 100) == 57) assign feedback = 19'h40269;
            else if((index % 100) == 58) assign feedback = 19'h4026C;
            else if((index % 100) == 59) assign feedback = 19'h4028E;
            else if((index % 100) == 60) assign feedback = 19'h40295;
            else if((index % 100) == 61) assign feedback = 19'h4029C;
            else if((index % 100) == 62) assign feedback = 19'h402A0;
            else if((index % 100) == 63) assign feedback = 19'h402A9;
            else if((index % 100) == 64) assign feedback = 19'h402AF;
            else if((index % 100) == 65) assign feedback = 19'h402B8;
            else if((index % 100) == 66) assign feedback = 19'h402BB;
            else if((index % 100) == 67) assign feedback = 19'h402D4;
            else if((index % 100) == 68) assign feedback = 19'h402DD;
            else if((index % 100) == 69) assign feedback = 19'h402E8;
            else if((index % 100) == 70) assign feedback = 19'h402EB;
            else if((index % 100) == 71) assign feedback = 19'h402EE;
            else if((index % 100) == 72) assign feedback = 19'h402F5;
            else if((index % 100) == 73) assign feedback = 19'h402FA;
            else if((index % 100) == 74) assign feedback = 19'h402FC;
            else if((index % 100) == 75) assign feedback = 19'h40304;
            else if((index % 100) == 76) assign feedback = 19'h40308;
            else if((index % 100) == 77) assign feedback = 19'h40319;
            else if((index % 100) == 78) assign feedback = 19'h40320;
            else if((index % 100) == 79) assign feedback = 19'h40325;
            else if((index % 100) == 80) assign feedback = 19'h40326;
            else if((index % 100) == 81) assign feedback = 19'h4032F;
            else if((index % 100) == 82) assign feedback = 19'h40332;
            else if((index % 100) == 83) assign feedback = 19'h40343;
            else if((index % 100) == 84) assign feedback = 19'h40345;
            else if((index % 100) == 85) assign feedback = 19'h4035E;
            else if((index % 100) == 86) assign feedback = 19'h40361;
            else if((index % 100) == 87) assign feedback = 19'h40368;
            else if((index % 100) == 88) assign feedback = 19'h40373;
            else if((index % 100) == 89) assign feedback = 19'h40376;
            else if((index % 100) == 90) assign feedback = 19'h4038A;
            else if((index % 100) == 91) assign feedback = 19'h4039D;
            else if((index % 100) == 92) assign feedback = 19'h403A2;
            else if((index % 100) == 93) assign feedback = 19'h403A4;
            else if((index % 100) == 94) assign feedback = 19'h403AB;
            else if((index % 100) == 95) assign feedback = 19'h403C2;
            else if((index % 100) == 96) assign feedback = 19'h403C8;
            else if((index % 100) == 97) assign feedback = 19'h403CE;
            else if((index % 100) == 98) assign feedback = 19'h403F7;
            else if((index % 100) == 99) assign feedback = 19'h403FE;
         end
      else if(width == 20)
         begin
            if((index % 100) == 0) assign feedback = 20'h80004;
            else if((index % 100) == 1) assign feedback = 20'h80029;
            else if((index % 100) == 2) assign feedback = 20'h80032;
            else if((index % 100) == 3) assign feedback = 20'h80034;
            else if((index % 100) == 4) assign feedback = 20'h8003D;
            else if((index % 100) == 5) assign feedback = 20'h80079;
            else if((index % 100) == 6) assign feedback = 20'h800B3;
            else if((index % 100) == 7) assign feedback = 20'h800B6;
            else if((index % 100) == 8) assign feedback = 20'h800BF;
            else if((index % 100) == 9) assign feedback = 20'h800C7;
            else if((index % 100) == 10) assign feedback = 20'h800DF;
            else if((index % 100) == 11) assign feedback = 20'h80111;
            else if((index % 100) == 12) assign feedback = 20'h80114;
            else if((index % 100) == 13) assign feedback = 20'h80118;
            else if((index % 100) == 14) assign feedback = 20'h8015C;
            else if((index % 100) == 15) assign feedback = 20'h80199;
            else if((index % 100) == 16) assign feedback = 20'h801A9;
            else if((index % 100) == 17) assign feedback = 20'h801AC;
            else if((index % 100) == 18) assign feedback = 20'h801B7;
            else if((index % 100) == 19) assign feedback = 20'h801E1;
            else if((index % 100) == 20) assign feedback = 20'h801FA;
            else if((index % 100) == 21) assign feedback = 20'h801FF;
            else if((index % 100) == 22) assign feedback = 20'h80211;
            else if((index % 100) == 23) assign feedback = 20'h80242;
            else if((index % 100) == 24) assign feedback = 20'h8024B;
            else if((index % 100) == 25) assign feedback = 20'h80260;
            else if((index % 100) == 26) assign feedback = 20'h80263;
            else if((index % 100) == 27) assign feedback = 20'h80266;
            else if((index % 100) == 28) assign feedback = 20'h80274;
            else if((index % 100) == 29) assign feedback = 20'h80284;
            else if((index % 100) == 30) assign feedback = 20'h80295;
            else if((index % 100) == 31) assign feedback = 20'h802CF;
            else if((index % 100) == 32) assign feedback = 20'h802F6;
            else if((index % 100) == 33) assign feedback = 20'h802F9;
            else if((index % 100) == 34) assign feedback = 20'h80302;
            else if((index % 100) == 35) assign feedback = 20'h80315;
            else if((index % 100) == 36) assign feedback = 20'h8031C;
            else if((index % 100) == 37) assign feedback = 20'h8032A;
            else if((index % 100) == 38) assign feedback = 20'h80338;
            else if((index % 100) == 39) assign feedback = 20'h8033D;
            else if((index % 100) == 40) assign feedback = 20'h8035B;
            else if((index % 100) == 41) assign feedback = 20'h8036E;
            else if((index % 100) == 42) assign feedback = 20'h80379;
            else if((index % 100) == 43) assign feedback = 20'h8038A;
            else if((index % 100) == 44) assign feedback = 20'h8039B;
            else if((index % 100) == 45) assign feedback = 20'h803A4;
            else if((index % 100) == 46) assign feedback = 20'h803BC;
            else if((index % 100) == 47) assign feedback = 20'h803EF;
            else if((index % 100) == 48) assign feedback = 20'h803FB;
            else if((index % 100) == 49) assign feedback = 20'h8040C;
            else if((index % 100) == 50) assign feedback = 20'h80414;
            else if((index % 100) == 51) assign feedback = 20'h8041B;
            else if((index % 100) == 52) assign feedback = 20'h80421;
            else if((index % 100) == 53) assign feedback = 20'h80448;
            else if((index % 100) == 54) assign feedback = 20'h8044D;
            else if((index % 100) == 55) assign feedback = 20'h80456;
            else if((index % 100) == 56) assign feedback = 20'h8045F;
            else if((index % 100) == 57) assign feedback = 20'h8048D;
            else if((index % 100) == 58) assign feedback = 20'h80499;
            else if((index % 100) == 59) assign feedback = 20'h8049C;
            else if((index % 100) == 60) assign feedback = 20'h804A6;
            else if((index % 100) == 61) assign feedback = 20'h804BD;
            else if((index % 100) == 62) assign feedback = 20'h804C6;
            else if((index % 100) == 63) assign feedback = 20'h804CC;
            else if((index % 100) == 64) assign feedback = 20'h804D7;
            else if((index % 100) == 65) assign feedback = 20'h804E7;
            else if((index % 100) == 66) assign feedback = 20'h804EE;
            else if((index % 100) == 67) assign feedback = 20'h804F0;
            else if((index % 100) == 68) assign feedback = 20'h80504;
            else if((index % 100) == 69) assign feedback = 20'h80513;
            else if((index % 100) == 70) assign feedback = 20'h8051A;
            else if((index % 100) == 71) assign feedback = 20'h80526;
            else if((index % 100) == 72) assign feedback = 20'h80529;
            else if((index % 100) == 73) assign feedback = 20'h80534;
            else if((index % 100) == 74) assign feedback = 20'h80543;
            else if((index % 100) == 75) assign feedback = 20'h8054A;
            else if((index % 100) == 76) assign feedback = 20'h80558;
            else if((index % 100) == 77) assign feedback = 20'h80568;
            else if((index % 100) == 78) assign feedback = 20'h8057A;
            else if((index % 100) == 79) assign feedback = 20'h805BC;
            else if((index % 100) == 80) assign feedback = 20'h805C1;
            else if((index % 100) == 81) assign feedback = 20'h805EA;
            else if((index % 100) == 82) assign feedback = 20'h805EC;
            else if((index % 100) == 83) assign feedback = 20'h80608;
            else if((index % 100) == 84) assign feedback = 20'h80637;
            else if((index % 100) == 85) assign feedback = 20'h8065B;
            else if((index % 100) == 86) assign feedback = 20'h8069D;
            else if((index % 100) == 87) assign feedback = 20'h8069E;
            else if((index % 100) == 88) assign feedback = 20'h806D0;
            else if((index % 100) == 89) assign feedback = 20'h80705;
            else if((index % 100) == 90) assign feedback = 20'h80718;
            else if((index % 100) == 91) assign feedback = 20'h80733;
            else if((index % 100) == 92) assign feedback = 20'h80735;
            else if((index % 100) == 93) assign feedback = 20'h80741;
            else if((index % 100) == 94) assign feedback = 20'h80753;
            else if((index % 100) == 95) assign feedback = 20'h80769;
            else if((index % 100) == 96) assign feedback = 20'h8076F;
            else if((index % 100) == 97) assign feedback = 20'h80799;
            else if((index % 100) == 98) assign feedback = 20'h807A5;
            else if((index % 100) == 99) assign feedback = 20'h807B8;
         end
      else if(width == 21)
         begin
            if((index % 100) == 0) assign feedback = 21'h100002;
            else if((index % 100) == 1) assign feedback = 21'h100013;
            else if((index % 100) == 2) assign feedback = 21'h10001F;
            else if((index % 100) == 3) assign feedback = 21'h100032;
            else if((index % 100) == 4) assign feedback = 21'h100037;
            else if((index % 100) == 5) assign feedback = 21'h10003D;
            else if((index % 100) == 6) assign feedback = 21'h10003E;
            else if((index % 100) == 7) assign feedback = 21'h100049;
            else if((index % 100) == 8) assign feedback = 21'h10005B;
            else if((index % 100) == 9) assign feedback = 21'h100083;
            else if((index % 100) == 10) assign feedback = 21'h10008F;
            else if((index % 100) == 11) assign feedback = 21'h10009D;
            else if((index % 100) == 12) assign feedback = 21'h1000A4;
            else if((index % 100) == 13) assign feedback = 21'h1000A7;
            else if((index % 100) == 14) assign feedback = 21'h1000B6;
            else if((index % 100) == 15) assign feedback = 21'h1000B9;
            else if((index % 100) == 16) assign feedback = 21'h1000C2;
            else if((index % 100) == 17) assign feedback = 21'h1000CB;
            else if((index % 100) == 18) assign feedback = 21'h1000CE;
            else if((index % 100) == 19) assign feedback = 21'h1000D3;
            else if((index % 100) == 20) assign feedback = 21'h1000D5;
            else if((index % 100) == 21) assign feedback = 21'h1000DA;
            else if((index % 100) == 22) assign feedback = 21'h1000DC;
            else if((index % 100) == 23) assign feedback = 21'h1000F1;
            else if((index % 100) == 24) assign feedback = 21'h1000F7;
            else if((index % 100) == 25) assign feedback = 21'h10010C;
            else if((index % 100) == 26) assign feedback = 21'h100112;
            else if((index % 100) == 27) assign feedback = 21'h10011B;
            else if((index % 100) == 28) assign feedback = 21'h10011E;
            else if((index % 100) == 29) assign feedback = 21'h10012D;
            else if((index % 100) == 30) assign feedback = 21'h100139;
            else if((index % 100) == 31) assign feedback = 21'h100156;
            else if((index % 100) == 32) assign feedback = 21'h100169;
            else if((index % 100) == 33) assign feedback = 21'h100184;
            else if((index % 100) == 34) assign feedback = 21'h10018D;
            else if((index % 100) == 35) assign feedback = 21'h1001A9;
            else if((index % 100) == 36) assign feedback = 21'h1001B1;
            else if((index % 100) == 37) assign feedback = 21'h1001BB;
            else if((index % 100) == 38) assign feedback = 21'h1001CF;
            else if((index % 100) == 39) assign feedback = 21'h1001D1;
            else if((index % 100) == 40) assign feedback = 21'h1001D7;
            else if((index % 100) == 41) assign feedback = 21'h1001DD;
            else if((index % 100) == 42) assign feedback = 21'h1001E2;
            else if((index % 100) == 43) assign feedback = 21'h1001EE;
            else if((index % 100) == 44) assign feedback = 21'h10020A;
            else if((index % 100) == 45) assign feedback = 21'h10020C;
            else if((index % 100) == 46) assign feedback = 21'h100211;
            else if((index % 100) == 47) assign feedback = 21'h100224;
            else if((index % 100) == 48) assign feedback = 21'h10022E;
            else if((index % 100) == 49) assign feedback = 21'h10023A;
            else if((index % 100) == 50) assign feedback = 21'h100248;
            else if((index % 100) == 51) assign feedback = 21'h10024B;
            else if((index % 100) == 52) assign feedback = 21'h100253;
            else if((index % 100) == 53) assign feedback = 21'h100272;
            else if((index % 100) == 54) assign feedback = 21'h100274;
            else if((index % 100) == 55) assign feedback = 21'h100277;
            else if((index % 100) == 56) assign feedback = 21'h10027E;
            else if((index % 100) == 57) assign feedback = 21'h100287;
            else if((index % 100) == 58) assign feedback = 21'h100295;
            else if((index % 100) == 59) assign feedback = 21'h1002AA;
            else if((index % 100) == 60) assign feedback = 21'h1002DB;
            else if((index % 100) == 61) assign feedback = 21'h1002EB;
            else if((index % 100) == 62) assign feedback = 21'h1002F0;
            else if((index % 100) == 63) assign feedback = 21'h1002F5;
            else if((index % 100) == 64) assign feedback = 21'h1002F6;
            else if((index % 100) == 65) assign feedback = 21'h100308;
            else if((index % 100) == 66) assign feedback = 21'h10031F;
            else if((index % 100) == 67) assign feedback = 21'h100329;
            else if((index % 100) == 68) assign feedback = 21'h100345;
            else if((index % 100) == 69) assign feedback = 21'h10035D;
            else if((index % 100) == 70) assign feedback = 21'h100361;
            else if((index % 100) == 71) assign feedback = 21'h10036B;
            else if((index % 100) == 72) assign feedback = 21'h100370;
            else if((index % 100) == 73) assign feedback = 21'h10037F;
            else if((index % 100) == 74) assign feedback = 21'h1003A1;
            else if((index % 100) == 75) assign feedback = 21'h1003AE;
            else if((index % 100) == 76) assign feedback = 21'h1003B5;
            else if((index % 100) == 77) assign feedback = 21'h1003BA;
            else if((index % 100) == 78) assign feedback = 21'h1003CB;
            else if((index % 100) == 79) assign feedback = 21'h1003D5;
            else if((index % 100) == 80) assign feedback = 21'h1003D9;
            else if((index % 100) == 81) assign feedback = 21'h1003E0;
            else if((index % 100) == 82) assign feedback = 21'h1003E6;
            else if((index % 100) == 83) assign feedback = 21'h1003E9;
            else if((index % 100) == 84) assign feedback = 21'h100406;
            else if((index % 100) == 85) assign feedback = 21'h100409;
            else if((index % 100) == 86) assign feedback = 21'h10040A;
            else if((index % 100) == 87) assign feedback = 21'h100427;
            else if((index % 100) == 88) assign feedback = 21'h100430;
            else if((index % 100) == 89) assign feedback = 21'h100441;
            else if((index % 100) == 90) assign feedback = 21'h100448;
            else if((index % 100) == 91) assign feedback = 21'h10044B;
            else if((index % 100) == 92) assign feedback = 21'h100455;
            else if((index % 100) == 93) assign feedback = 21'h10045C;
            else if((index % 100) == 94) assign feedback = 21'h10046F;
            else if((index % 100) == 95) assign feedback = 21'h100478;
            else if((index % 100) == 96) assign feedback = 21'h10047D;
            else if((index % 100) == 97) assign feedback = 21'h10049A;
            else if((index % 100) == 98) assign feedback = 21'h1004AC;
            else if((index % 100) == 99) assign feedback = 21'h1004B2;
         end
      else if(width == 22)
         begin
            if((index % 100) == 0) assign feedback = 22'h200001;
            else if((index % 100) == 1) assign feedback = 22'h20001C;
            else if((index % 100) == 2) assign feedback = 22'h20005E;
            else if((index % 100) == 3) assign feedback = 22'h200061;
            else if((index % 100) == 4) assign feedback = 22'h200094;
            else if((index % 100) == 5) assign feedback = 22'h2000B0;
            else if((index % 100) == 6) assign feedback = 22'h2000B9;
            else if((index % 100) == 7) assign feedback = 22'h2000C7;
            else if((index % 100) == 8) assign feedback = 22'h2000D9;
            else if((index % 100) == 9) assign feedback = 22'h2000F8;
            else if((index % 100) == 10) assign feedback = 22'h200111;
            else if((index % 100) == 11) assign feedback = 22'h200133;
            else if((index % 100) == 12) assign feedback = 22'h200156;
            else if((index % 100) == 13) assign feedback = 22'h20015A;
            else if((index % 100) == 14) assign feedback = 22'h200182;
            else if((index % 100) == 15) assign feedback = 22'h200188;
            else if((index % 100) == 16) assign feedback = 22'h2001A5;
            else if((index % 100) == 17) assign feedback = 22'h2001B4;
            else if((index % 100) == 18) assign feedback = 22'h2001C0;
            else if((index % 100) == 19) assign feedback = 22'h2001DB;
            else if((index % 100) == 20) assign feedback = 22'h2001E7;
            else if((index % 100) == 21) assign feedback = 22'h2001EB;
            else if((index % 100) == 22) assign feedback = 22'h2001ED;
            else if((index % 100) == 23) assign feedback = 22'h200209;
            else if((index % 100) == 24) assign feedback = 22'h200239;
            else if((index % 100) == 25) assign feedback = 22'h200244;
            else if((index % 100) == 26) assign feedback = 22'h200272;
            else if((index % 100) == 27) assign feedback = 22'h200287;
            else if((index % 100) == 28) assign feedback = 22'h20028D;
            else if((index % 100) == 29) assign feedback = 22'h20029F;
            else if((index % 100) == 30) assign feedback = 22'h2002A3;
            else if((index % 100) == 31) assign feedback = 22'h2002BD;
            else if((index % 100) == 32) assign feedback = 22'h2002C3;
            else if((index % 100) == 33) assign feedback = 22'h2002C6;
            else if((index % 100) == 34) assign feedback = 22'h2002CC;
            else if((index % 100) == 35) assign feedback = 22'h2002DD;
            else if((index % 100) == 36) assign feedback = 22'h20030B;
            else if((index % 100) == 37) assign feedback = 22'h20030D;
            else if((index % 100) == 38) assign feedback = 22'h200332;
            else if((index % 100) == 39) assign feedback = 22'h200345;
            else if((index % 100) == 40) assign feedback = 22'h200358;
            else if((index % 100) == 41) assign feedback = 22'h200361;
            else if((index % 100) == 42) assign feedback = 22'h20036D;
            else if((index % 100) == 43) assign feedback = 22'h200398;
            else if((index % 100) == 44) assign feedback = 22'h2003B5;
            else if((index % 100) == 45) assign feedback = 22'h2003BF;
            else if((index % 100) == 46) assign feedback = 22'h2003C2;
            else if((index % 100) == 47) assign feedback = 22'h2003E3;
            else if((index % 100) == 48) assign feedback = 22'h2003EC;
            else if((index % 100) == 49) assign feedback = 22'h2003FD;
            else if((index % 100) == 50) assign feedback = 22'h200403;
            else if((index % 100) == 51) assign feedback = 22'h200414;
            else if((index % 100) == 52) assign feedback = 22'h200427;
            else if((index % 100) == 53) assign feedback = 22'h200433;
            else if((index % 100) == 54) assign feedback = 22'h20044B;
            else if((index % 100) == 55) assign feedback = 22'h200459;
            else if((index % 100) == 56) assign feedback = 22'h200460;
            else if((index % 100) == 57) assign feedback = 22'h200463;
            else if((index % 100) == 58) assign feedback = 22'h200481;
            else if((index % 100) == 59) assign feedback = 22'h20049F;
            else if((index % 100) == 60) assign feedback = 22'h2004BE;
            else if((index % 100) == 61) assign feedback = 22'h2004C6;
            else if((index % 100) == 62) assign feedback = 22'h2004D7;
            else if((index % 100) == 63) assign feedback = 22'h2004DD;
            else if((index % 100) == 64) assign feedback = 22'h2004E1;
            else if((index % 100) == 65) assign feedback = 22'h2004E2;
            else if((index % 100) == 66) assign feedback = 22'h2004ED;
            else if((index % 100) == 67) assign feedback = 22'h2004FA;
            else if((index % 100) == 68) assign feedback = 22'h200515;
            else if((index % 100) == 69) assign feedback = 22'h20051C;
            else if((index % 100) == 70) assign feedback = 22'h20053E;
            else if((index % 100) == 71) assign feedback = 22'h20054A;
            else if((index % 100) == 72) assign feedback = 22'h20054F;
            else if((index % 100) == 73) assign feedback = 22'h20056E;
            else if((index % 100) == 74) assign feedback = 22'h200575;
            else if((index % 100) == 75) assign feedback = 22'h200576;
            else if((index % 100) == 76) assign feedback = 22'h20057C;
            else if((index % 100) == 77) assign feedback = 22'h200589;
            else if((index % 100) == 78) assign feedback = 22'h2005A4;
            else if((index % 100) == 79) assign feedback = 22'h2005AD;
            else if((index % 100) == 80) assign feedback = 22'h2005B3;
            else if((index % 100) == 81) assign feedback = 22'h2005B6;
            else if((index % 100) == 82) assign feedback = 22'h2005BA;
            else if((index % 100) == 83) assign feedback = 22'h2005BF;
            else if((index % 100) == 84) assign feedback = 22'h2005EC;
            else if((index % 100) == 85) assign feedback = 22'h2005EF;
            else if((index % 100) == 86) assign feedback = 22'h200616;
            else if((index % 100) == 87) assign feedback = 22'h200623;
            else if((index % 100) == 88) assign feedback = 22'h200634;
            else if((index % 100) == 89) assign feedback = 22'h20064A;
            else if((index % 100) == 90) assign feedback = 22'h20064C;
            else if((index % 100) == 91) assign feedback = 22'h20064F;
            else if((index % 100) == 92) assign feedback = 22'h200651;
            else if((index % 100) == 93) assign feedback = 22'h200667;
            else if((index % 100) == 94) assign feedback = 22'h20066B;
            else if((index % 100) == 95) assign feedback = 22'h200685;
            else if((index % 100) == 96) assign feedback = 22'h200697;
            else if((index % 100) == 97) assign feedback = 22'h20069B;
            else if((index % 100) == 98) assign feedback = 22'h20069E;
            else if((index % 100) == 99) assign feedback = 22'h2006A8;
         end
      else if(width == 23)
         begin
            if((index % 100) == 0) assign feedback = 23'h400010;
            else if((index % 100) == 1) assign feedback = 23'h400015;
            else if((index % 100) == 2) assign feedback = 23'h400016;
            else if((index % 100) == 3) assign feedback = 23'h400019;
            else if((index % 100) == 4) assign feedback = 23'h40001F;
            else if((index % 100) == 5) assign feedback = 23'h400026;
            else if((index % 100) == 6) assign feedback = 23'h400032;
            else if((index % 100) == 7) assign feedback = 23'h40003B;
            else if((index % 100) == 8) assign feedback = 23'h400043;
            else if((index % 100) == 9) assign feedback = 23'h400045;
            else if((index % 100) == 10) assign feedback = 23'h40004C;
            else if((index % 100) == 11) assign feedback = 23'h400051;
            else if((index % 100) == 12) assign feedback = 23'h40005E;
            else if((index % 100) == 13) assign feedback = 23'h400062;
            else if((index % 100) == 14) assign feedback = 23'h400079;
            else if((index % 100) == 15) assign feedback = 23'h40007C;
            else if((index % 100) == 16) assign feedback = 23'h400097;
            else if((index % 100) == 17) assign feedback = 23'h40009D;
            else if((index % 100) == 18) assign feedback = 23'h4000AD;
            else if((index % 100) == 19) assign feedback = 23'h4000B0;
            else if((index % 100) == 20) assign feedback = 23'h4000B3;
            else if((index % 100) == 21) assign feedback = 23'h4000C1;
            else if((index % 100) == 22) assign feedback = 23'h4000C4;
            else if((index % 100) == 23) assign feedback = 23'h4000FB;
            else if((index % 100) == 24) assign feedback = 23'h400100;
            else if((index % 100) == 25) assign feedback = 23'h40010F;
            else if((index % 100) == 26) assign feedback = 23'h400112;
            else if((index % 100) == 27) assign feedback = 23'h400124;
            else if((index % 100) == 28) assign feedback = 23'h400127;
            else if((index % 100) == 29) assign feedback = 23'h40012B;
            else if((index % 100) == 30) assign feedback = 23'h40012D;
            else if((index % 100) == 31) assign feedback = 23'h400136;
            else if((index % 100) == 32) assign feedback = 23'h40013C;
            else if((index % 100) == 33) assign feedback = 23'h400147;
            else if((index % 100) == 34) assign feedback = 23'h400148;
            else if((index % 100) == 35) assign feedback = 23'h40015C;
            else if((index % 100) == 36) assign feedback = 23'h40016F;
            else if((index % 100) == 37) assign feedback = 23'h400177;
            else if((index % 100) == 38) assign feedback = 23'h400181;
            else if((index % 100) == 39) assign feedback = 23'h400193;
            else if((index % 100) == 40) assign feedback = 23'h400196;
            else if((index % 100) == 41) assign feedback = 23'h4001A0;
            else if((index % 100) == 42) assign feedback = 23'h4001B2;
            else if((index % 100) == 43) assign feedback = 23'h4001D1;
            else if((index % 100) == 44) assign feedback = 23'h4001D2;
            else if((index % 100) == 45) assign feedback = 23'h4001D8;
            else if((index % 100) == 46) assign feedback = 23'h4001DE;
            else if((index % 100) == 47) assign feedback = 23'h4001F6;
            else if((index % 100) == 48) assign feedback = 23'h400206;
            else if((index % 100) == 49) assign feedback = 23'h400214;
            else if((index % 100) == 50) assign feedback = 23'h400228;
            else if((index % 100) == 51) assign feedback = 23'h400247;
            else if((index % 100) == 52) assign feedback = 23'h400260;
            else if((index % 100) == 53) assign feedback = 23'h40026F;
            else if((index % 100) == 54) assign feedback = 23'h400293;
            else if((index % 100) == 55) assign feedback = 23'h400295;
            else if((index % 100) == 56) assign feedback = 23'h4002A0;
            else if((index % 100) == 57) assign feedback = 23'h4002B7;
            else if((index % 100) == 58) assign feedback = 23'h4002D2;
            else if((index % 100) == 59) assign feedback = 23'h4002D4;
            else if((index % 100) == 60) assign feedback = 23'h4002E2;
            else if((index % 100) == 61) assign feedback = 23'h4002F0;
            else if((index % 100) == 62) assign feedback = 23'h400308;
            else if((index % 100) == 63) assign feedback = 23'h40030E;
            else if((index % 100) == 64) assign feedback = 23'h40032F;
            else if((index % 100) == 65) assign feedback = 23'h400331;
            else if((index % 100) == 66) assign feedback = 23'h400340;
            else if((index % 100) == 67) assign feedback = 23'h40035D;
            else if((index % 100) == 68) assign feedback = 23'h400362;
            else if((index % 100) == 69) assign feedback = 23'h40036D;
            else if((index % 100) == 70) assign feedback = 23'h40036E;
            else if((index % 100) == 71) assign feedback = 23'h400376;
            else if((index % 100) == 72) assign feedback = 23'h400379;
            else if((index % 100) == 73) assign feedback = 23'h400389;
            else if((index % 100) == 74) assign feedback = 23'h40038A;
            else if((index % 100) == 75) assign feedback = 23'h400391;
            else if((index % 100) == 76) assign feedback = 23'h40039B;
            else if((index % 100) == 77) assign feedback = 23'h4003BF;
            else if((index % 100) == 78) assign feedback = 23'h4003D0;
            else if((index % 100) == 79) assign feedback = 23'h4003DA;
            else if((index % 100) == 80) assign feedback = 23'h4003EF;
            else if((index % 100) == 81) assign feedback = 23'h4003F2;
            else if((index % 100) == 82) assign feedback = 23'h4003FB;
            else if((index % 100) == 83) assign feedback = 23'h4003FD;
            else if((index % 100) == 84) assign feedback = 23'h40041D;
            else if((index % 100) == 85) assign feedback = 23'h40041E;
            else if((index % 100) == 86) assign feedback = 23'h40042D;
            else if((index % 100) == 87) assign feedback = 23'h40043F;
            else if((index % 100) == 88) assign feedback = 23'h400444;
            else if((index % 100) == 89) assign feedback = 23'h40044D;
            else if((index % 100) == 90) assign feedback = 23'h400455;
            else if((index % 100) == 91) assign feedback = 23'h400456;
            else if((index % 100) == 92) assign feedback = 23'h400460;
            else if((index % 100) == 93) assign feedback = 23'h400463;
            else if((index % 100) == 94) assign feedback = 23'h40046A;
            else if((index % 100) == 95) assign feedback = 23'h400484;
            else if((index % 100) == 96) assign feedback = 23'h400490;
            else if((index % 100) == 97) assign feedback = 23'h40049C;
            else if((index % 100) == 98) assign feedback = 23'h4004AA;
            else if((index % 100) == 99) assign feedback = 23'h4004B2;
         end
      else if(width == 24)
         begin
            if((index % 100) == 0) assign feedback = 24'h80000D;
            else if((index % 100) == 1) assign feedback = 24'h800043;
            else if((index % 100) == 2) assign feedback = 24'h800058;
            else if((index % 100) == 3) assign feedback = 24'h80006D;
            else if((index % 100) == 4) assign feedback = 24'h80007A;
            else if((index % 100) == 5) assign feedback = 24'h800092;
            else if((index % 100) == 6) assign feedback = 24'h8000BF;
            else if((index % 100) == 7) assign feedback = 24'h8000DA;
            else if((index % 100) == 8) assign feedback = 24'h8000E5;
            else if((index % 100) == 9) assign feedback = 24'h800112;
            else if((index % 100) == 10) assign feedback = 24'h800128;
            else if((index % 100) == 11) assign feedback = 24'h80012B;
            else if((index % 100) == 12) assign feedback = 24'h800136;
            else if((index % 100) == 13) assign feedback = 24'h8001B1;
            else if((index % 100) == 14) assign feedback = 24'h8001B4;
            else if((index % 100) == 15) assign feedback = 24'h8001D7;
            else if((index % 100) == 16) assign feedback = 24'h8001E1;
            else if((index % 100) == 17) assign feedback = 24'h8001E7;
            else if((index % 100) == 18) assign feedback = 24'h8001F9;
            else if((index % 100) == 19) assign feedback = 24'h80020C;
            else if((index % 100) == 20) assign feedback = 24'h800221;
            else if((index % 100) == 21) assign feedback = 24'h800224;
            else if((index % 100) == 22) assign feedback = 24'h8002BD;
            else if((index % 100) == 23) assign feedback = 24'h800329;
            else if((index % 100) == 24) assign feedback = 24'h800345;
            else if((index % 100) == 25) assign feedback = 24'h80035E;
            else if((index % 100) == 26) assign feedback = 24'h8003A7;
            else if((index % 100) == 27) assign feedback = 24'h8003A8;
            else if((index % 100) == 28) assign feedback = 24'h8003C7;
            else if((index % 100) == 29) assign feedback = 24'h800412;
            else if((index % 100) == 30) assign feedback = 24'h80041B;
            else if((index % 100) == 31) assign feedback = 24'h800422;
            else if((index % 100) == 32) assign feedback = 24'h80042B;
            else if((index % 100) == 33) assign feedback = 24'h80044E;
            else if((index % 100) == 34) assign feedback = 24'h800453;
            else if((index % 100) == 35) assign feedback = 24'h80047E;
            else if((index % 100) == 36) assign feedback = 24'h800481;
            else if((index % 100) == 37) assign feedback = 24'h8004DE;
            else if((index % 100) == 38) assign feedback = 24'h8004ED;
            else if((index % 100) == 39) assign feedback = 24'h8004F6;
            else if((index % 100) == 40) assign feedback = 24'h800507;
            else if((index % 100) == 41) assign feedback = 24'h800520;
            else if((index % 100) == 42) assign feedback = 24'h800523;
            else if((index % 100) == 43) assign feedback = 24'h80053D;
            else if((index % 100) == 44) assign feedback = 24'h80055D;
            else if((index % 100) == 45) assign feedback = 24'h800579;
            else if((index % 100) == 46) assign feedback = 24'h800580;
            else if((index % 100) == 47) assign feedback = 24'h80058F;
            else if((index % 100) == 48) assign feedback = 24'h800594;
            else if((index % 100) == 49) assign feedback = 24'h80059B;
            else if((index % 100) == 50) assign feedback = 24'h8005A2;
            else if((index % 100) == 51) assign feedback = 24'h8005A4;
            else if((index % 100) == 52) assign feedback = 24'h8005A8;
            else if((index % 100) == 53) assign feedback = 24'h8005BA;
            else if((index % 100) == 54) assign feedback = 24'h8005D6;
            else if((index % 100) == 55) assign feedback = 24'h8005EA;
            else if((index % 100) == 56) assign feedback = 24'h800602;
            else if((index % 100) == 57) assign feedback = 24'h800613;
            else if((index % 100) == 58) assign feedback = 24'h80066E;
            else if((index % 100) == 59) assign feedback = 24'h80067F;
            else if((index % 100) == 60) assign feedback = 24'h80069B;
            else if((index % 100) == 61) assign feedback = 24'h8006B5;
            else if((index % 100) == 62) assign feedback = 24'h8006E6;
            else if((index % 100) == 63) assign feedback = 24'h8006E9;
            else if((index % 100) == 64) assign feedback = 24'h8006EF;
            else if((index % 100) == 65) assign feedback = 24'h8006F4;
            else if((index % 100) == 66) assign feedback = 24'h80070A;
            else if((index % 100) == 67) assign feedback = 24'h800730;
            else if((index % 100) == 68) assign feedback = 24'h800759;
            else if((index % 100) == 69) assign feedback = 24'h80075F;
            else if((index % 100) == 70) assign feedback = 24'h800795;
            else if((index % 100) == 71) assign feedback = 24'h8007BE;
            else if((index % 100) == 72) assign feedback = 24'h8007DE;
            else if((index % 100) == 73) assign feedback = 24'h8007E4;
            else if((index % 100) == 74) assign feedback = 24'h800806;
            else if((index % 100) == 75) assign feedback = 24'h800817;
            else if((index % 100) == 76) assign feedback = 24'h800853;
            else if((index % 100) == 77) assign feedback = 24'h800863;
            else if((index % 100) == 78) assign feedback = 24'h8008A6;
            else if((index % 100) == 79) assign feedback = 24'h8008D1;
            else if((index % 100) == 80) assign feedback = 24'h8008D7;
            else if((index % 100) == 81) assign feedback = 24'h8008E7;
            else if((index % 100) == 82) assign feedback = 24'h8008F3;
            else if((index % 100) == 83) assign feedback = 24'h8008FC;
            else if((index % 100) == 84) assign feedback = 24'h80090B;
            else if((index % 100) == 85) assign feedback = 24'h800916;
            else if((index % 100) == 86) assign feedback = 24'h80093B;
            else if((index % 100) == 87) assign feedback = 24'h800973;
            else if((index % 100) == 88) assign feedback = 24'h8009F8;
            else if((index % 100) == 89) assign feedback = 24'h8009FE;
            else if((index % 100) == 90) assign feedback = 24'h800A23;
            else if((index % 100) == 91) assign feedback = 24'h800A3E;
            else if((index % 100) == 92) assign feedback = 24'h800AA1;
            else if((index % 100) == 93) assign feedback = 24'h800AA7;
            else if((index % 100) == 94) assign feedback = 24'h800AAB;
            else if((index % 100) == 95) assign feedback = 24'h800AC4;
            else if((index % 100) == 96) assign feedback = 24'h800AD5;
            else if((index % 100) == 97) assign feedback = 24'h800B35;
            else if((index % 100) == 98) assign feedback = 24'h800B4D;
            else if((index % 100) == 99) assign feedback = 24'h800B87;
         end
      else if(width == 25)
         begin
            if((index % 100) == 0) assign feedback = 25'h1000004;
            else if((index % 100) == 1) assign feedback = 25'h1000007;
            else if((index % 100) == 2) assign feedback = 25'h1000016;
            else if((index % 100) == 3) assign feedback = 25'h1000040;
            else if((index % 100) == 4) assign feedback = 25'h1000049;
            else if((index % 100) == 5) assign feedback = 25'h1000062;
            else if((index % 100) == 6) assign feedback = 25'h100007F;
            else if((index % 100) == 7) assign feedback = 25'h1000086;
            else if((index % 100) == 8) assign feedback = 25'h100009E;
            else if((index % 100) == 9) assign feedback = 25'h10000A2;
            else if((index % 100) == 10) assign feedback = 25'h10000B9;
            else if((index % 100) == 11) assign feedback = 25'h10000CB;
            else if((index % 100) == 12) assign feedback = 25'h10000D0;
            else if((index % 100) == 13) assign feedback = 25'h10000D6;
            else if((index % 100) == 14) assign feedback = 25'h10000DC;
            else if((index % 100) == 15) assign feedback = 25'h10000E9;
            else if((index % 100) == 16) assign feedback = 25'h10000EF;
            else if((index % 100) == 17) assign feedback = 25'h10000F4;
            else if((index % 100) == 18) assign feedback = 25'h100010A;
            else if((index % 100) == 19) assign feedback = 25'h1000111;
            else if((index % 100) == 20) assign feedback = 25'h1000118;
            else if((index % 100) == 21) assign feedback = 25'h1000144;
            else if((index % 100) == 22) assign feedback = 25'h1000160;
            else if((index % 100) == 23) assign feedback = 25'h1000165;
            else if((index % 100) == 24) assign feedback = 25'h100016F;
            else if((index % 100) == 25) assign feedback = 25'h1000172;
            else if((index % 100) == 26) assign feedback = 25'h100017D;
            else if((index % 100) == 27) assign feedback = 25'h1000182;
            else if((index % 100) == 28) assign feedback = 25'h100018B;
            else if((index % 100) == 29) assign feedback = 25'h1000190;
            else if((index % 100) == 30) assign feedback = 25'h100019C;
            else if((index % 100) == 31) assign feedback = 25'h10001A5;
            else if((index % 100) == 32) assign feedback = 25'h10001A6;
            else if((index % 100) == 33) assign feedback = 25'h10001AF;
            else if((index % 100) == 34) assign feedback = 25'h10001B7;
            else if((index % 100) == 35) assign feedback = 25'h10001E2;
            else if((index % 100) == 36) assign feedback = 25'h10001F5;
            else if((index % 100) == 37) assign feedback = 25'h10001FC;
            else if((index % 100) == 38) assign feedback = 25'h1000205;
            else if((index % 100) == 39) assign feedback = 25'h1000206;
            else if((index % 100) == 40) assign feedback = 25'h1000239;
            else if((index % 100) == 41) assign feedback = 25'h100025F;
            else if((index % 100) == 42) assign feedback = 25'h100026A;
            else if((index % 100) == 43) assign feedback = 25'h1000272;
            else if((index % 100) == 44) assign feedback = 25'h100027B;
            else if((index % 100) == 45) assign feedback = 25'h100027E;
            else if((index % 100) == 46) assign feedback = 25'h1000287;
            else if((index % 100) == 47) assign feedback = 25'h1000290;
            else if((index % 100) == 48) assign feedback = 25'h1000296;
            else if((index % 100) == 49) assign feedback = 25'h100029F;
            else if((index % 100) == 50) assign feedback = 25'h10002A3;
            else if((index % 100) == 51) assign feedback = 25'h10002B4;
            else if((index % 100) == 52) assign feedback = 25'h10002B8;
            else if((index % 100) == 53) assign feedback = 25'h10002D8;
            else if((index % 100) == 54) assign feedback = 25'h10002E7;
            else if((index % 100) == 55) assign feedback = 25'h10002EB;
            else if((index % 100) == 56) assign feedback = 25'h10002F3;
            else if((index % 100) == 57) assign feedback = 25'h1000310;
            else if((index % 100) == 58) assign feedback = 25'h1000319;
            else if((index % 100) == 59) assign feedback = 25'h1000320;
            else if((index % 100) == 60) assign feedback = 25'h100032F;
            else if((index % 100) == 61) assign feedback = 25'h1000334;
            else if((index % 100) == 62) assign feedback = 25'h100033D;
            else if((index % 100) == 63) assign feedback = 25'h1000349;
            else if((index % 100) == 64) assign feedback = 25'h100035B;
            else if((index % 100) == 65) assign feedback = 25'h1000361;
            else if((index % 100) == 66) assign feedback = 25'h1000376;
            else if((index % 100) == 67) assign feedback = 25'h100037C;
            else if((index % 100) == 68) assign feedback = 25'h1000386;
            else if((index % 100) == 69) assign feedback = 25'h1000392;
            else if((index % 100) == 70) assign feedback = 25'h1000398;
            else if((index % 100) == 71) assign feedback = 25'h100039B;
            else if((index % 100) == 72) assign feedback = 25'h100039D;
            else if((index % 100) == 73) assign feedback = 25'h10003C8;
            else if((index % 100) == 74) assign feedback = 25'h10003CE;
            else if((index % 100) == 75) assign feedback = 25'h10003DA;
            else if((index % 100) == 76) assign feedback = 25'h10003DC;
            else if((index % 100) == 77) assign feedback = 25'h10003E5;
            else if((index % 100) == 78) assign feedback = 25'h10003EA;
            else if((index % 100) == 79) assign feedback = 25'h10003F1;
            else if((index % 100) == 80) assign feedback = 25'h10003FD;
            else if((index % 100) == 81) assign feedback = 25'h100042B;
            else if((index % 100) == 82) assign feedback = 25'h100042E;
            else if((index % 100) == 83) assign feedback = 25'h100043A;
            else if((index % 100) == 84) assign feedback = 25'h1000444;
            else if((index % 100) == 85) assign feedback = 25'h100044E;
            else if((index % 100) == 86) assign feedback = 25'h1000469;
            else if((index % 100) == 87) assign feedback = 25'h100046A;
            else if((index % 100) == 88) assign feedback = 25'h1000478;
            else if((index % 100) == 89) assign feedback = 25'h100047B;
            else if((index % 100) == 90) assign feedback = 25'h100048D;
            else if((index % 100) == 91) assign feedback = 25'h100048E;
            else if((index % 100) == 92) assign feedback = 25'h1000493;
            else if((index % 100) == 93) assign feedback = 25'h1000495;
            else if((index % 100) == 94) assign feedback = 25'h10004A0;
            else if((index % 100) == 95) assign feedback = 25'h10004B1;
            else if((index % 100) == 96) assign feedback = 25'h10004B7;
            else if((index % 100) == 97) assign feedback = 25'h10004C9;
            else if((index % 100) == 98) assign feedback = 25'h10004EB;
            else if((index % 100) == 99) assign feedback = 25'h10004F3;
         end
      else if(width == 26)
         begin
            if((index % 100) == 0) assign feedback = 26'h2000023;
            else if((index % 100) == 1) assign feedback = 26'h2000026;
            else if((index % 100) == 2) assign feedback = 26'h2000058;
            else if((index % 100) == 3) assign feedback = 26'h2000070;
            else if((index % 100) == 4) assign feedback = 26'h200007A;
            else if((index % 100) == 5) assign feedback = 26'h200008C;
            else if((index % 100) == 6) assign feedback = 26'h200009D;
            else if((index % 100) == 7) assign feedback = 26'h20000B6;
            else if((index % 100) == 8) assign feedback = 26'h20000BF;
            else if((index % 100) == 9) assign feedback = 26'h20000C1;
            else if((index % 100) == 10) assign feedback = 26'h20000C4;
            else if((index % 100) == 11) assign feedback = 26'h20000DF;
            else if((index % 100) == 12) assign feedback = 26'h20000F1;
            else if((index % 100) == 13) assign feedback = 26'h2000109;
            else if((index % 100) == 14) assign feedback = 26'h200011D;
            else if((index % 100) == 15) assign feedback = 26'h2000122;
            else if((index % 100) == 16) assign feedback = 26'h2000139;
            else if((index % 100) == 17) assign feedback = 26'h2000142;
            else if((index % 100) == 18) assign feedback = 26'h200014E;
            else if((index % 100) == 19) assign feedback = 26'h2000155;
            else if((index % 100) == 20) assign feedback = 26'h200015C;
            else if((index % 100) == 21) assign feedback = 26'h2000178;
            else if((index % 100) == 22) assign feedback = 26'h200017D;
            else if((index % 100) == 23) assign feedback = 26'h20001A0;
            else if((index % 100) == 24) assign feedback = 26'h20001A5;
            else if((index % 100) == 25) assign feedback = 26'h20001DB;
            else if((index % 100) == 26) assign feedback = 26'h20001E4;
            else if((index % 100) == 27) assign feedback = 26'h20001FC;
            else if((index % 100) == 28) assign feedback = 26'h2000214;
            else if((index % 100) == 29) assign feedback = 26'h200021D;
            else if((index % 100) == 30) assign feedback = 26'h2000244;
            else if((index % 100) == 31) assign feedback = 26'h200024B;
            else if((index % 100) == 32) assign feedback = 26'h200024D;
            else if((index % 100) == 33) assign feedback = 26'h2000250;
            else if((index % 100) == 34) assign feedback = 26'h2000274;
            else if((index % 100) == 35) assign feedback = 26'h200028E;
            else if((index % 100) == 36) assign feedback = 26'h20002BE;
            else if((index % 100) == 37) assign feedback = 26'h20002C5;
            else if((index % 100) == 38) assign feedback = 26'h20002DB;
            else if((index % 100) == 39) assign feedback = 26'h20002E2;
            else if((index % 100) == 40) assign feedback = 26'h2000323;
            else if((index % 100) == 41) assign feedback = 26'h2000331;
            else if((index % 100) == 42) assign feedback = 26'h200033D;
            else if((index % 100) == 43) assign feedback = 26'h2000346;
            else if((index % 100) == 44) assign feedback = 26'h200034A;
            else if((index % 100) == 45) assign feedback = 26'h2000376;
            else if((index % 100) == 46) assign feedback = 26'h200037F;
            else if((index % 100) == 47) assign feedback = 26'h2000383;
            else if((index % 100) == 48) assign feedback = 26'h2000385;
            else if((index % 100) == 49) assign feedback = 26'h200038C;
            else if((index % 100) == 50) assign feedback = 26'h2000398;
            else if((index % 100) == 51) assign feedback = 26'h200039B;
            else if((index % 100) == 52) assign feedback = 26'h200039E;
            else if((index % 100) == 53) assign feedback = 26'h20003A7;
            else if((index % 100) == 54) assign feedback = 26'h20003D6;
            else if((index % 100) == 55) assign feedback = 26'h2000414;
            else if((index % 100) == 56) assign feedback = 26'h200041B;
            else if((index % 100) == 57) assign feedback = 26'h2000421;
            else if((index % 100) == 58) assign feedback = 26'h200042D;
            else if((index % 100) == 59) assign feedback = 26'h200045F;
            else if((index % 100) == 60) assign feedback = 26'h2000460;
            else if((index % 100) == 61) assign feedback = 26'h2000472;
            else if((index % 100) == 62) assign feedback = 26'h2000477;
            else if((index % 100) == 63) assign feedback = 26'h2000484;
            else if((index % 100) == 64) assign feedback = 26'h2000487;
            else if((index % 100) == 65) assign feedback = 26'h2000495;
            else if((index % 100) == 66) assign feedback = 26'h20004CC;
            else if((index % 100) == 67) assign feedback = 26'h20004D8;
            else if((index % 100) == 68) assign feedback = 26'h20004DE;
            else if((index % 100) == 69) assign feedback = 26'h200051A;
            else if((index % 100) == 70) assign feedback = 26'h200053E;
            else if((index % 100) == 71) assign feedback = 26'h200055B;
            else if((index % 100) == 72) assign feedback = 26'h200057A;
            else if((index % 100) == 73) assign feedback = 26'h2000580;
            else if((index % 100) == 74) assign feedback = 26'h2000589;
            else if((index % 100) == 75) assign feedback = 26'h2000592;
            else if((index % 100) == 76) assign feedback = 26'h20005A7;
            else if((index % 100) == 77) assign feedback = 26'h20005BC;
            else if((index % 100) == 78) assign feedback = 26'h20005BF;
            else if((index % 100) == 79) assign feedback = 26'h20005C2;
            else if((index % 100) == 80) assign feedback = 26'h20005D5;
            else if((index % 100) == 81) assign feedback = 26'h20005DA;
            else if((index % 100) == 82) assign feedback = 26'h20005E3;
            else if((index % 100) == 83) assign feedback = 26'h20005F1;
            else if((index % 100) == 84) assign feedback = 26'h2000607;
            else if((index % 100) == 85) assign feedback = 26'h2000608;
            else if((index % 100) == 86) assign feedback = 26'h200062C;
            else if((index % 100) == 87) assign feedback = 26'h2000637;
            else if((index % 100) == 88) assign feedback = 26'h2000645;
            else if((index % 100) == 89) assign feedback = 26'h200065B;
            else if((index % 100) == 90) assign feedback = 26'h2000679;
            else if((index % 100) == 91) assign feedback = 26'h200068F;
            else if((index % 100) == 92) assign feedback = 26'h20006B9;
            else if((index % 100) == 93) assign feedback = 26'h20006CD;
            else if((index % 100) == 94) assign feedback = 26'h20006D5;
            else if((index % 100) == 95) assign feedback = 26'h20006E3;
            else if((index % 100) == 96) assign feedback = 26'h20006F4;
            else if((index % 100) == 97) assign feedback = 26'h2000700;
            else if((index % 100) == 98) assign feedback = 26'h2000709;
            else if((index % 100) == 99) assign feedback = 26'h200072D;
         end
      else if(width == 27)
         begin
            if((index % 100) == 0) assign feedback = 27'h4000013;
            else if((index % 100) == 1) assign feedback = 27'h4000068;
            else if((index % 100) == 2) assign feedback = 27'h4000073;
            else if((index % 100) == 3) assign feedback = 27'h4000075;
            else if((index % 100) == 4) assign feedback = 27'h4000094;
            else if((index % 100) == 5) assign feedback = 27'h4000098;
            else if((index % 100) == 6) assign feedback = 27'h40000AE;
            else if((index % 100) == 7) assign feedback = 27'h40000B6;
            else if((index % 100) == 8) assign feedback = 27'h40000BC;
            else if((index % 100) == 9) assign feedback = 27'h40000C1;
            else if((index % 100) == 10) assign feedback = 27'h40000F1;
            else if((index % 100) == 11) assign feedback = 27'h4000112;
            else if((index % 100) == 12) assign feedback = 27'h4000114;
            else if((index % 100) == 13) assign feedback = 27'h400011B;
            else if((index % 100) == 14) assign feedback = 27'h4000128;
            else if((index % 100) == 15) assign feedback = 27'h4000144;
            else if((index % 100) == 16) assign feedback = 27'h4000182;
            else if((index % 100) == 17) assign feedback = 27'h40001AA;
            else if((index % 100) == 18) assign feedback = 27'h40001B4;
            else if((index % 100) == 19) assign feedback = 27'h40001BD;
            else if((index % 100) == 20) assign feedback = 27'h40001D1;
            else if((index % 100) == 21) assign feedback = 27'h40001D4;
            else if((index % 100) == 22) assign feedback = 27'h40001E7;
            else if((index % 100) == 23) assign feedback = 27'h4000203;
            else if((index % 100) == 24) assign feedback = 27'h4000218;
            else if((index % 100) == 25) assign feedback = 27'h4000227;
            else if((index % 100) == 26) assign feedback = 27'h400022D;
            else if((index % 100) == 27) assign feedback = 27'h400022E;
            else if((index % 100) == 28) assign feedback = 27'h4000242;
            else if((index % 100) == 29) assign feedback = 27'h400024D;
            else if((index % 100) == 30) assign feedback = 27'h400025A;
            else if((index % 100) == 31) assign feedback = 27'h4000277;
            else if((index % 100) == 32) assign feedback = 27'h4000290;
            else if((index % 100) == 33) assign feedback = 27'h40002A5;
            else if((index % 100) == 34) assign feedback = 27'h40002AA;
            else if((index % 100) == 35) assign feedback = 27'h40002B7;
            else if((index % 100) == 36) assign feedback = 27'h40002C0;
            else if((index % 100) == 37) assign feedback = 27'h40002D2;
            else if((index % 100) == 38) assign feedback = 27'h40002D8;
            else if((index % 100) == 39) assign feedback = 27'h40002F0;
            else if((index % 100) == 40) assign feedback = 27'h40002F5;
            else if((index % 100) == 41) assign feedback = 27'h40002FC;
            else if((index % 100) == 42) assign feedback = 27'h400031A;
            else if((index % 100) == 43) assign feedback = 27'h400031C;
            else if((index % 100) == 44) assign feedback = 27'h400032C;
            else if((index % 100) == 45) assign feedback = 27'h4000340;
            else if((index % 100) == 46) assign feedback = 27'h400034C;
            else if((index % 100) == 47) assign feedback = 27'h4000354;
            else if((index % 100) == 48) assign feedback = 27'h400035D;
            else if((index % 100) == 49) assign feedback = 27'h400039E;
            else if((index % 100) == 50) assign feedback = 27'h40003A7;
            else if((index % 100) == 51) assign feedback = 27'h40003AB;
            else if((index % 100) == 52) assign feedback = 27'h40003B3;
            else if((index % 100) == 53) assign feedback = 27'h40003B5;
            else if((index % 100) == 54) assign feedback = 27'h40003B9;
            else if((index % 100) == 55) assign feedback = 27'h40003DF;
            else if((index % 100) == 56) assign feedback = 27'h40003E3;
            else if((index % 100) == 57) assign feedback = 27'h40003F4;
            else if((index % 100) == 58) assign feedback = 27'h400040F;
            else if((index % 100) == 59) assign feedback = 27'h400042B;
            else if((index % 100) == 60) assign feedback = 27'h4000436;
            else if((index % 100) == 61) assign feedback = 27'h4000453;
            else if((index % 100) == 62) assign feedback = 27'h4000471;
            else if((index % 100) == 63) assign feedback = 27'h4000474;
            else if((index % 100) == 64) assign feedback = 27'h400048D;
            else if((index % 100) == 65) assign feedback = 27'h4000499;
            else if((index % 100) == 66) assign feedback = 27'h40004A6;
            else if((index % 100) == 67) assign feedback = 27'h40004B2;
            else if((index % 100) == 68) assign feedback = 27'h40004BD;
            else if((index % 100) == 69) assign feedback = 27'h40004D1;
            else if((index % 100) == 70) assign feedback = 27'h40004DB;
            else if((index % 100) == 71) assign feedback = 27'h40004E7;
            else if((index % 100) == 72) assign feedback = 27'h40004ED;
            else if((index % 100) == 73) assign feedback = 27'h40004F5;
            else if((index % 100) == 74) assign feedback = 27'h4000507;
            else if((index % 100) == 75) assign feedback = 27'h400050E;
            else if((index % 100) == 76) assign feedback = 27'h400052A;
            else if((index % 100) == 77) assign feedback = 27'h4000534;
            else if((index % 100) == 78) assign feedback = 27'h4000545;
            else if((index % 100) == 79) assign feedback = 27'h400054C;
            else if((index % 100) == 80) assign feedback = 27'h4000551;
            else if((index % 100) == 81) assign feedback = 27'h4000562;
            else if((index % 100) == 82) assign feedback = 27'h400056E;
            else if((index % 100) == 83) assign feedback = 27'h4000597;
            else if((index % 100) == 84) assign feedback = 27'h400059E;
            else if((index % 100) == 85) assign feedback = 27'h40005A4;
            else if((index % 100) == 86) assign feedback = 27'h40005BF;
            else if((index % 100) == 87) assign feedback = 27'h40005D3;
            else if((index % 100) == 88) assign feedback = 27'h40005D6;
            else if((index % 100) == 89) assign feedback = 27'h40005E9;
            else if((index % 100) == 90) assign feedback = 27'h40005EC;
            else if((index % 100) == 91) assign feedback = 27'h40005FB;
            else if((index % 100) == 92) assign feedback = 27'h4000607;
            else if((index % 100) == 93) assign feedback = 27'h400062F;
            else if((index % 100) == 94) assign feedback = 27'h4000649;
            else if((index % 100) == 95) assign feedback = 27'h4000652;
            else if((index % 100) == 96) assign feedback = 27'h4000670;
            else if((index % 100) == 97) assign feedback = 27'h400067C;
            else if((index % 100) == 98) assign feedback = 27'h4000680;
            else if((index % 100) == 99) assign feedback = 27'h40006AE;
         end
      else if(width == 28)
         begin
            if((index % 100) == 0) assign feedback = 28'h8000004;
            else if((index % 100) == 1) assign feedback = 28'h8000029;
            else if((index % 100) == 2) assign feedback = 28'h800003B;
            else if((index % 100) == 3) assign feedback = 28'h8000070;
            else if((index % 100) == 4) assign feedback = 28'h80000B3;
            else if((index % 100) == 5) assign feedback = 28'h80000B9;
            else if((index % 100) == 6) assign feedback = 28'h80000EF;
            else if((index % 100) == 7) assign feedback = 28'h8000100;
            else if((index % 100) == 8) assign feedback = 28'h8000111;
            else if((index % 100) == 9) assign feedback = 28'h8000159;
            else if((index % 100) == 10) assign feedback = 28'h800016C;
            else if((index % 100) == 11) assign feedback = 28'h8000190;
            else if((index % 100) == 12) assign feedback = 28'h800019C;
            else if((index % 100) == 13) assign feedback = 28'h80001AC;
            else if((index % 100) == 14) assign feedback = 28'h80001B8;
            else if((index % 100) == 15) assign feedback = 28'h80001D8;
            else if((index % 100) == 16) assign feedback = 28'h8000205;
            else if((index % 100) == 17) assign feedback = 28'h8000214;
            else if((index % 100) == 18) assign feedback = 28'h8000217;
            else if((index % 100) == 19) assign feedback = 28'h8000256;
            else if((index % 100) == 20) assign feedback = 28'h800025A;
            else if((index % 100) == 21) assign feedback = 28'h800027E;
            else if((index % 100) == 22) assign feedback = 28'h8000296;
            else if((index % 100) == 23) assign feedback = 28'h80002E1;
            else if((index % 100) == 24) assign feedback = 28'h80002EB;
            else if((index % 100) == 25) assign feedback = 28'h80002F5;
            else if((index % 100) == 26) assign feedback = 28'h8000308;
            else if((index % 100) == 27) assign feedback = 28'h800031F;
            else if((index % 100) == 28) assign feedback = 28'h8000334;
            else if((index % 100) == 29) assign feedback = 28'h800033E;
            else if((index % 100) == 30) assign feedback = 28'h8000358;
            else if((index % 100) == 31) assign feedback = 28'h800035B;
            else if((index % 100) == 32) assign feedback = 28'h800037F;
            else if((index % 100) == 33) assign feedback = 28'h8000380;
            else if((index % 100) == 34) assign feedback = 28'h8000386;
            else if((index % 100) == 35) assign feedback = 28'h80003C8;
            else if((index % 100) == 36) assign feedback = 28'h80003CB;
            else if((index % 100) == 37) assign feedback = 28'h80003E6;
            else if((index % 100) == 38) assign feedback = 28'h800043A;
            else if((index % 100) == 39) assign feedback = 28'h8000444;
            else if((index % 100) == 40) assign feedback = 28'h800044B;
            else if((index % 100) == 41) assign feedback = 28'h8000456;
            else if((index % 100) == 42) assign feedback = 28'h800047D;
            else if((index % 100) == 43) assign feedback = 28'h800048D;
            else if((index % 100) == 44) assign feedback = 28'h800049A;
            else if((index % 100) == 45) assign feedback = 28'h80004B2;
            else if((index % 100) == 46) assign feedback = 28'h80004BB;
            else if((index % 100) == 47) assign feedback = 28'h80004D2;
            else if((index % 100) == 48) assign feedback = 28'h80004D7;
            else if((index % 100) == 49) assign feedback = 28'h80004E8;
            else if((index % 100) == 50) assign feedback = 28'h800050E;
            else if((index % 100) == 51) assign feedback = 28'h8000554;
            else if((index % 100) == 52) assign feedback = 28'h8000564;
            else if((index % 100) == 53) assign feedback = 28'h800056B;
            else if((index % 100) == 54) assign feedback = 28'h8000579;
            else if((index % 100) == 55) assign feedback = 28'h800057C;
            else if((index % 100) == 56) assign feedback = 28'h8000597;
            else if((index % 100) == 57) assign feedback = 28'h80005AD;
            else if((index % 100) == 58) assign feedback = 28'h80005C1;
            else if((index % 100) == 59) assign feedback = 28'h80005C2;
            else if((index % 100) == 60) assign feedback = 28'h80005E6;
            else if((index % 100) == 61) assign feedback = 28'h80005F7;
            else if((index % 100) == 62) assign feedback = 28'h8000604;
            else if((index % 100) == 63) assign feedback = 28'h8000662;
            else if((index % 100) == 64) assign feedback = 28'h8000668;
            else if((index % 100) == 65) assign feedback = 28'h800068F;
            else if((index % 100) == 66) assign feedback = 28'h800069D;
            else if((index % 100) == 67) assign feedback = 28'h80006BA;
            else if((index % 100) == 68) assign feedback = 28'h80006CE;
            else if((index % 100) == 69) assign feedback = 28'h80006FB;
            else if((index % 100) == 70) assign feedback = 28'h800070F;
            else if((index % 100) == 71) assign feedback = 28'h8000724;
            else if((index % 100) == 72) assign feedback = 28'h8000727;
            else if((index % 100) == 73) assign feedback = 28'h8000735;
            else if((index % 100) == 74) assign feedback = 28'h80007A5;
            else if((index % 100) == 75) assign feedback = 28'h80007A9;
            else if((index % 100) == 76) assign feedback = 28'h80007AF;
            else if((index % 100) == 77) assign feedback = 28'h80007DB;
            else if((index % 100) == 78) assign feedback = 28'h80007F3;
            else if((index % 100) == 79) assign feedback = 28'h80007F6;
            else if((index % 100) == 80) assign feedback = 28'h80007FF;
            else if((index % 100) == 81) assign feedback = 28'h8000803;
            else if((index % 100) == 82) assign feedback = 28'h800082D;
            else if((index % 100) == 83) assign feedback = 28'h8000835;
            else if((index % 100) == 84) assign feedback = 28'h8000836;
            else if((index % 100) == 85) assign feedback = 28'h8000853;
            else if((index % 100) == 86) assign feedback = 28'h8000893;
            else if((index % 100) == 87) assign feedback = 28'h80008E2;
            else if((index % 100) == 88) assign feedback = 28'h8000907;
            else if((index % 100) == 89) assign feedback = 28'h800090E;
            else if((index % 100) == 90) assign feedback = 28'h800092C;
            else if((index % 100) == 91) assign feedback = 28'h8000932;
            else if((index % 100) == 92) assign feedback = 28'h8000949;
            else if((index % 100) == 93) assign feedback = 28'h8000961;
            else if((index % 100) == 94) assign feedback = 28'h8000964;
            else if((index % 100) == 95) assign feedback = 28'h8000979;
            else if((index % 100) == 96) assign feedback = 28'h8000991;
            else if((index % 100) == 97) assign feedback = 28'h80009AE;
            else if((index % 100) == 98) assign feedback = 28'h80009DC;
            else if((index % 100) == 99) assign feedback = 28'h80009E3;
         end
      else if(width == 29)
         begin
            if((index % 100) == 0) assign feedback = 29'h10000002;
            else if((index % 100) == 1) assign feedback = 29'h1000000B;
            else if((index % 100) == 2) assign feedback = 29'h1000000E;
            else if((index % 100) == 3) assign feedback = 29'h10000046;
            else if((index % 100) == 4) assign feedback = 29'h10000061;
            else if((index % 100) == 5) assign feedback = 29'h1000007C;
            else if((index % 100) == 6) assign feedback = 29'h1000008C;
            else if((index % 100) == 7) assign feedback = 29'h1000009D;
            else if((index % 100) == 8) assign feedback = 29'h1000009E;
            else if((index % 100) == 9) assign feedback = 29'h100000B9;
            else if((index % 100) == 10) assign feedback = 29'h100000C4;
            else if((index % 100) == 11) assign feedback = 29'h100000C8;
            else if((index % 100) == 12) assign feedback = 29'h100000D5;
            else if((index % 100) == 13) assign feedback = 29'h100000DF;
            else if((index % 100) == 14) assign feedback = 29'h10000103;
            else if((index % 100) == 15) assign feedback = 29'h1000010A;
            else if((index % 100) == 16) assign feedback = 29'h10000130;
            else if((index % 100) == 17) assign feedback = 29'h10000139;
            else if((index % 100) == 18) assign feedback = 29'h10000147;
            else if((index % 100) == 19) assign feedback = 29'h10000182;
            else if((index % 100) == 20) assign feedback = 29'h100001A5;
            else if((index % 100) == 21) assign feedback = 29'h100001A9;
            else if((index % 100) == 22) assign feedback = 29'h100001B2;
            else if((index % 100) == 23) assign feedback = 29'h100001BB;
            else if((index % 100) == 24) assign feedback = 29'h100001BE;
            else if((index % 100) == 25) assign feedback = 29'h100001CA;
            else if((index % 100) == 26) assign feedback = 29'h100001DE;
            else if((index % 100) == 27) assign feedback = 29'h100001FA;
            else if((index % 100) == 28) assign feedback = 29'h10000206;
            else if((index % 100) == 29) assign feedback = 29'h10000211;
            else if((index % 100) == 30) assign feedback = 29'h10000218;
            else if((index % 100) == 31) assign feedback = 29'h10000221;
            else if((index % 100) == 32) assign feedback = 29'h1000022E;
            else if((index % 100) == 33) assign feedback = 29'h10000235;
            else if((index % 100) == 34) assign feedback = 29'h10000239;
            else if((index % 100) == 35) assign feedback = 29'h1000023C;
            else if((index % 100) == 36) assign feedback = 29'h1000024B;
            else if((index % 100) == 37) assign feedback = 29'h1000024D;
            else if((index % 100) == 38) assign feedback = 29'h10000256;
            else if((index % 100) == 39) assign feedback = 29'h10000260;
            else if((index % 100) == 40) assign feedback = 29'h1000026F;
            else if((index % 100) == 41) assign feedback = 29'h1000027B;
            else if((index % 100) == 42) assign feedback = 29'h1000029A;
            else if((index % 100) == 43) assign feedback = 29'h1000029F;
            else if((index % 100) == 44) assign feedback = 29'h100002A0;
            else if((index % 100) == 45) assign feedback = 29'h100002A5;
            else if((index % 100) == 46) assign feedback = 29'h100002A9;
            else if((index % 100) == 47) assign feedback = 29'h100002B8;
            else if((index % 100) == 48) assign feedback = 29'h100002C5;
            else if((index % 100) == 49) assign feedback = 29'h100002D7;
            else if((index % 100) == 50) assign feedback = 29'h100002DD;
            else if((index % 100) == 51) assign feedback = 29'h100002E2;
            else if((index % 100) == 52) assign feedback = 29'h100002EB;
            else if((index % 100) == 53) assign feedback = 29'h100002F3;
            else if((index % 100) == 54) assign feedback = 29'h10000308;
            else if((index % 100) == 55) assign feedback = 29'h10000310;
            else if((index % 100) == 56) assign feedback = 29'h1000031A;
            else if((index % 100) == 57) assign feedback = 29'h10000331;
            else if((index % 100) == 58) assign feedback = 29'h10000337;
            else if((index % 100) == 59) assign feedback = 29'h10000340;
            else if((index % 100) == 60) assign feedback = 29'h10000349;
            else if((index % 100) == 61) assign feedback = 29'h10000352;
            else if((index % 100) == 62) assign feedback = 29'h10000370;
            else if((index % 100) == 63) assign feedback = 29'h10000375;
            else if((index % 100) == 64) assign feedback = 29'h10000385;
            else if((index % 100) == 65) assign feedback = 29'h10000389;
            else if((index % 100) == 66) assign feedback = 29'h1000038A;
            else if((index % 100) == 67) assign feedback = 29'h1000038C;
            else if((index % 100) == 68) assign feedback = 29'h10000398;
            else if((index % 100) == 69) assign feedback = 29'h100003A8;
            else if((index % 100) == 70) assign feedback = 29'h100003C1;
            else if((index % 100) == 71) assign feedback = 29'h100003C2;
            else if((index % 100) == 72) assign feedback = 29'h100003D3;
            else if((index % 100) == 73) assign feedback = 29'h100003D6;
            else if((index % 100) == 74) assign feedback = 29'h100003E6;
            else if((index % 100) == 75) assign feedback = 29'h100003FD;
            else if((index % 100) == 76) assign feedback = 29'h1000041E;
            else if((index % 100) == 77) assign feedback = 29'h10000422;
            else if((index % 100) == 78) assign feedback = 29'h1000042D;
            else if((index % 100) == 79) assign feedback = 29'h10000447;
            else if((index % 100) == 80) assign feedback = 29'h10000455;
            else if((index % 100) == 81) assign feedback = 29'h10000460;
            else if((index % 100) == 82) assign feedback = 29'h1000046C;
            else if((index % 100) == 83) assign feedback = 29'h10000471;
            else if((index % 100) == 84) assign feedback = 29'h100004A9;
            else if((index % 100) == 85) assign feedback = 29'h100004B1;
            else if((index % 100) == 86) assign feedback = 29'h100004B2;
            else if((index % 100) == 87) assign feedback = 29'h100004B4;
            else if((index % 100) == 88) assign feedback = 29'h100004BB;
            else if((index % 100) == 89) assign feedback = 29'h100004C6;
            else if((index % 100) == 90) assign feedback = 29'h100004F3;
            else if((index % 100) == 91) assign feedback = 29'h10000502;
            else if((index % 100) == 92) assign feedback = 29'h10000508;
            else if((index % 100) == 93) assign feedback = 29'h1000051F;
            else if((index % 100) == 94) assign feedback = 29'h10000557;
            else if((index % 100) == 95) assign feedback = 29'h1000055B;
            else if((index % 100) == 96) assign feedback = 29'h1000055E;
            else if((index % 100) == 97) assign feedback = 29'h10000564;
            else if((index % 100) == 98) assign feedback = 29'h10000576;
            else if((index % 100) == 99) assign feedback = 29'h10000583;
         end
      else if(width == 30)
         begin
            if((index % 100) == 0) assign feedback = 30'h20000029;
            else if((index % 100) == 1) assign feedback = 30'h20000057;
            else if((index % 100) == 2) assign feedback = 30'h2000005E;
            else if((index % 100) == 3) assign feedback = 30'h20000089;
            else if((index % 100) == 4) assign feedback = 30'h200000A4;
            else if((index % 100) == 5) assign feedback = 30'h200000EC;
            else if((index % 100) == 6) assign feedback = 30'h2000011E;
            else if((index % 100) == 7) assign feedback = 30'h20000148;
            else if((index % 100) == 8) assign feedback = 30'h2000014E;
            else if((index % 100) == 9) assign feedback = 30'h20000160;
            else if((index % 100) == 10) assign feedback = 30'h20000172;
            else if((index % 100) == 11) assign feedback = 30'h2000017B;
            else if((index % 100) == 12) assign feedback = 30'h2000018B;
            else if((index % 100) == 13) assign feedback = 30'h200001E7;
            else if((index % 100) == 14) assign feedback = 30'h200001EB;
            else if((index % 100) == 15) assign feedback = 30'h20000241;
            else if((index % 100) == 16) assign feedback = 30'h20000244;
            else if((index % 100) == 17) assign feedback = 30'h2000027B;
            else if((index % 100) == 18) assign feedback = 30'h2000027D;
            else if((index % 100) == 19) assign feedback = 30'h200002AC;
            else if((index % 100) == 20) assign feedback = 30'h2000031A;
            else if((index % 100) == 21) assign feedback = 30'h20000332;
            else if((index % 100) == 22) assign feedback = 30'h20000354;
            else if((index % 100) == 23) assign feedback = 30'h20000357;
            else if((index % 100) == 24) assign feedback = 30'h2000039E;
            else if((index % 100) == 25) assign feedback = 30'h200003AB;
            else if((index % 100) == 26) assign feedback = 30'h200003B9;
            else if((index % 100) == 27) assign feedback = 30'h2000041D;
            else if((index % 100) == 28) assign feedback = 30'h20000427;
            else if((index % 100) == 29) assign feedback = 30'h20000439;
            else if((index % 100) == 30) assign feedback = 30'h2000044E;
            else if((index % 100) == 31) assign feedback = 30'h2000046C;
            else if((index % 100) == 32) assign feedback = 30'h200004A5;
            else if((index % 100) == 33) assign feedback = 30'h200004BE;
            else if((index % 100) == 34) assign feedback = 30'h200004C5;
            else if((index % 100) == 35) assign feedback = 30'h200004C9;
            else if((index % 100) == 36) assign feedback = 30'h200004E1;
            else if((index % 100) == 37) assign feedback = 30'h200004E4;
            else if((index % 100) == 38) assign feedback = 30'h200004EE;
            else if((index % 100) == 39) assign feedback = 30'h2000054C;
            else if((index % 100) == 40) assign feedback = 30'h20000567;
            else if((index % 100) == 41) assign feedback = 30'h20000597;
            else if((index % 100) == 42) assign feedback = 30'h200005BA;
            else if((index % 100) == 43) assign feedback = 30'h20000602;
            else if((index % 100) == 44) assign feedback = 30'h20000619;
            else if((index % 100) == 45) assign feedback = 30'h2000061C;
            else if((index % 100) == 46) assign feedback = 30'h2000064A;
            else if((index % 100) == 47) assign feedback = 30'h2000065B;
            else if((index % 100) == 48) assign feedback = 30'h2000065D;
            else if((index % 100) == 49) assign feedback = 30'h20000679;
            else if((index % 100) == 50) assign feedback = 30'h200006CB;
            else if((index % 100) == 51) assign feedback = 30'h200006D3;
            else if((index % 100) == 52) assign feedback = 30'h20000705;
            else if((index % 100) == 53) assign feedback = 30'h20000735;
            else if((index % 100) == 54) assign feedback = 30'h20000759;
            else if((index % 100) == 55) assign feedback = 30'h200007D2;
            else if((index % 100) == 56) assign feedback = 30'h200007DD;
            else if((index % 100) == 57) assign feedback = 30'h200007EB;
            else if((index % 100) == 58) assign feedback = 30'h2000080F;
            else if((index % 100) == 59) assign feedback = 30'h20000841;
            else if((index % 100) == 60) assign feedback = 30'h20000847;
            else if((index % 100) == 61) assign feedback = 30'h2000084E;
            else if((index % 100) == 62) assign feedback = 30'h2000088D;
            else if((index % 100) == 63) assign feedback = 30'h200008B4;
            else if((index % 100) == 64) assign feedback = 30'h200008C3;
            else if((index % 100) == 65) assign feedback = 30'h200008DD;
            else if((index % 100) == 66) assign feedback = 30'h200008EB;
            else if((index % 100) == 67) assign feedback = 30'h20000910;
            else if((index % 100) == 68) assign feedback = 30'h2000093D;
            else if((index % 100) == 69) assign feedback = 30'h20000951;
            else if((index % 100) == 70) assign feedback = 30'h2000096E;
            else if((index % 100) == 71) assign feedback = 30'h20000998;
            else if((index % 100) == 72) assign feedback = 30'h2000099B;
            else if((index % 100) == 73) assign feedback = 30'h200009AD;
            else if((index % 100) == 74) assign feedback = 30'h200009C2;
            else if((index % 100) == 75) assign feedback = 30'h200009C8;
            else if((index % 100) == 76) assign feedback = 30'h200009D5;
            else if((index % 100) == 77) assign feedback = 30'h20000A45;
            else if((index % 100) == 78) assign feedback = 30'h20000A46;
            else if((index % 100) == 79) assign feedback = 30'h20000A9D;
            else if((index % 100) == 80) assign feedback = 30'h20000AE0;
            else if((index % 100) == 81) assign feedback = 30'h20000AE9;
            else if((index % 100) == 82) assign feedback = 30'h20000B03;
            else if((index % 100) == 83) assign feedback = 30'h20000B09;
            else if((index % 100) == 84) assign feedback = 30'h20000B18;
            else if((index % 100) == 85) assign feedback = 30'h20000B53;
            else if((index % 100) == 86) assign feedback = 30'h20000B72;
            else if((index % 100) == 87) assign feedback = 30'h20000B7D;
            else if((index % 100) == 88) assign feedback = 30'h20000B8E;
            else if((index % 100) == 89) assign feedback = 30'h20000BA3;
            else if((index % 100) == 90) assign feedback = 30'h20000BB8;
            else if((index % 100) == 91) assign feedback = 30'h20000BBE;
            else if((index % 100) == 92) assign feedback = 30'h20000BCA;
            else if((index % 100) == 93) assign feedback = 30'h20000BD1;
            else if((index % 100) == 94) assign feedback = 30'h20000C04;
            else if((index % 100) == 95) assign feedback = 30'h20000C10;
            else if((index % 100) == 96) assign feedback = 30'h20000C23;
            else if((index % 100) == 97) assign feedback = 30'h20000C34;
            else if((index % 100) == 98) assign feedback = 30'h20000C86;
            else if((index % 100) == 99) assign feedback = 30'h20000C92;
         end
      else if(width == 31)
         begin
            if((index % 100) == 0) assign feedback = 31'h40000004;
            else if((index % 100) == 1) assign feedback = 31'h40000007;
            else if((index % 100) == 2) assign feedback = 31'h40000016;
            else if((index % 100) == 3) assign feedback = 31'h4000001A;
            else if((index % 100) == 4) assign feedback = 31'h40000020;
            else if((index % 100) == 5) assign feedback = 31'h40000023;
            else if((index % 100) == 6) assign feedback = 31'h4000002A;
            else if((index % 100) == 7) assign feedback = 31'h40000040;
            else if((index % 100) == 8) assign feedback = 31'h40000045;
            else if((index % 100) == 9) assign feedback = 31'h40000054;
            else if((index % 100) == 10) assign feedback = 31'h4000005D;
            else if((index % 100) == 11) assign feedback = 31'h4000007F;
            else if((index % 100) == 12) assign feedback = 31'h4000008F;
            else if((index % 100) == 13) assign feedback = 31'h40000097;
            else if((index % 100) == 14) assign feedback = 31'h400000A2;
            else if((index % 100) == 15) assign feedback = 31'h400000AE;
            else if((index % 100) == 16) assign feedback = 31'h400000B0;
            else if((index % 100) == 17) assign feedback = 31'h400000B5;
            else if((index % 100) == 18) assign feedback = 31'h400000D0;
            else if((index % 100) == 19) assign feedback = 31'h400000D6;
            else if((index % 100) == 20) assign feedback = 31'h400000E3;
            else if((index % 100) == 21) assign feedback = 31'h40000105;
            else if((index % 100) == 22) assign feedback = 31'h40000111;
            else if((index % 100) == 23) assign feedback = 31'h40000118;
            else if((index % 100) == 24) assign feedback = 31'h4000013C;
            else if((index % 100) == 25) assign feedback = 31'h40000159;
            else if((index % 100) == 26) assign feedback = 31'h40000169;
            else if((index % 100) == 27) assign feedback = 31'h4000016F;
            else if((index % 100) == 28) assign feedback = 31'h4000017B;
            else if((index % 100) == 29) assign feedback = 31'h40000188;
            else if((index % 100) == 30) assign feedback = 31'h4000018E;
            else if((index % 100) == 31) assign feedback = 31'h40000193;
            else if((index % 100) == 32) assign feedback = 31'h400001BD;
            else if((index % 100) == 33) assign feedback = 31'h400001C9;
            else if((index % 100) == 34) assign feedback = 31'h400001ED;
            else if((index % 100) == 35) assign feedback = 31'h40000217;
            else if((index % 100) == 36) assign feedback = 31'h40000230;
            else if((index % 100) == 37) assign feedback = 31'h40000233;
            else if((index % 100) == 38) assign feedback = 31'h40000255;
            else if((index % 100) == 39) assign feedback = 31'h40000265;
            else if((index % 100) == 40) assign feedback = 31'h4000026A;
            else if((index % 100) == 41) assign feedback = 31'h40000272;
            else if((index % 100) == 42) assign feedback = 31'h40000278;
            else if((index % 100) == 43) assign feedback = 31'h4000028D;
            else if((index % 100) == 44) assign feedback = 31'h4000029C;
            else if((index % 100) == 45) assign feedback = 31'h4000029F;
            else if((index % 100) == 46) assign feedback = 31'h400002B8;
            else if((index % 100) == 47) assign feedback = 31'h400002C3;
            else if((index % 100) == 48) assign feedback = 31'h400002C6;
            else if((index % 100) == 49) assign feedback = 31'h400002E8;
            else if((index % 100) == 50) assign feedback = 31'h400002F3;
            else if((index % 100) == 51) assign feedback = 31'h400002FA;
            else if((index % 100) == 52) assign feedback = 31'h40000301;
            else if((index % 100) == 53) assign feedback = 31'h40000326;
            else if((index % 100) == 54) assign feedback = 31'h4000033B;
            else if((index % 100) == 55) assign feedback = 31'h4000034A;
            else if((index % 100) == 56) assign feedback = 31'h4000034C;
            else if((index % 100) == 57) assign feedback = 31'h4000037F;
            else if((index % 100) == 58) assign feedback = 31'h4000038F;
            else if((index % 100) == 59) assign feedback = 31'h40000394;
            else if((index % 100) == 60) assign feedback = 31'h4000039D;
            else if((index % 100) == 61) assign feedback = 31'h400003A4;
            else if((index % 100) == 62) assign feedback = 31'h400003B6;
            else if((index % 100) == 63) assign feedback = 31'h400003BF;
            else if((index % 100) == 64) assign feedback = 31'h400003C1;
            else if((index % 100) == 65) assign feedback = 31'h400003CB;
            else if((index % 100) == 66) assign feedback = 31'h400003DA;
            else if((index % 100) == 67) assign feedback = 31'h400003DC;
            else if((index % 100) == 68) assign feedback = 31'h400003EA;
            else if((index % 100) == 69) assign feedback = 31'h400003FE;
            else if((index % 100) == 70) assign feedback = 31'h40000403;
            else if((index % 100) == 71) assign feedback = 31'h4000040C;
            else if((index % 100) == 72) assign feedback = 31'h40000459;
            else if((index % 100) == 73) assign feedback = 31'h4000045C;
            else if((index % 100) == 74) assign feedback = 31'h4000045F;
            else if((index % 100) == 75) assign feedback = 31'h4000046A;
            else if((index % 100) == 76) assign feedback = 31'h40000474;
            else if((index % 100) == 77) assign feedback = 31'h4000047B;
            else if((index % 100) == 78) assign feedback = 31'h40000481;
            else if((index % 100) == 79) assign feedback = 31'h4000048D;
            else if((index % 100) == 80) assign feedback = 31'h40000493;
            else if((index % 100) == 81) assign feedback = 31'h400004B8;
            else if((index % 100) == 82) assign feedback = 31'h400004DE;
            else if((index % 100) == 83) assign feedback = 31'h400004ED;
            else if((index % 100) == 84) assign feedback = 31'h40000501;
            else if((index % 100) == 85) assign feedback = 31'h40000513;
            else if((index % 100) == 86) assign feedback = 31'h40000525;
            else if((index % 100) == 87) assign feedback = 31'h4000052F;
            else if((index % 100) == 88) assign feedback = 31'h40000534;
            else if((index % 100) == 89) assign feedback = 31'h40000538;
            else if((index % 100) == 90) assign feedback = 31'h4000053E;
            else if((index % 100) == 91) assign feedback = 31'h40000540;
            else if((index % 100) == 92) assign feedback = 31'h40000549;
            else if((index % 100) == 93) assign feedback = 31'h4000054F;
            else if((index % 100) == 94) assign feedback = 31'h4000055D;
            else if((index % 100) == 95) assign feedback = 31'h40000567;
            else if((index % 100) == 96) assign feedback = 31'h4000056B;
            else if((index % 100) == 97) assign feedback = 31'h40000576;
            else if((index % 100) == 98) assign feedback = 31'h40000585;
            else if((index % 100) == 99) assign feedback = 31'h400005B6;
         end
      else if(width == 32)
         begin
            if((index % 100) == 0) assign feedback = 32'h80000057;
            else if((index % 100) == 1) assign feedback = 32'h80000062;
            else if((index % 100) == 2) assign feedback = 32'h8000007A;
            else if((index % 100) == 3) assign feedback = 32'h80000092;
            else if((index % 100) == 4) assign feedback = 32'h800000B9;
            else if((index % 100) == 5) assign feedback = 32'h800000BA;
            else if((index % 100) == 6) assign feedback = 32'h80000106;
            else if((index % 100) == 7) assign feedback = 32'h80000114;
            else if((index % 100) == 8) assign feedback = 32'h8000012D;
            else if((index % 100) == 9) assign feedback = 32'h8000014E;
            else if((index % 100) == 10) assign feedback = 32'h8000016C;
            else if((index % 100) == 11) assign feedback = 32'h8000019F;
            else if((index % 100) == 12) assign feedback = 32'h800001A6;
            else if((index % 100) == 13) assign feedback = 32'h800001F3;
            else if((index % 100) == 14) assign feedback = 32'h8000020F;
            else if((index % 100) == 15) assign feedback = 32'h800002CC;
            else if((index % 100) == 16) assign feedback = 32'h80000349;
            else if((index % 100) == 17) assign feedback = 32'h80000370;
            else if((index % 100) == 18) assign feedback = 32'h80000375;
            else if((index % 100) == 19) assign feedback = 32'h80000392;
            else if((index % 100) == 20) assign feedback = 32'h80000398;
            else if((index % 100) == 21) assign feedback = 32'h800003BF;
            else if((index % 100) == 22) assign feedback = 32'h800003D6;
            else if((index % 100) == 23) assign feedback = 32'h800003DF;
            else if((index % 100) == 24) assign feedback = 32'h800003E9;
            else if((index % 100) == 25) assign feedback = 32'h80000412;
            else if((index % 100) == 26) assign feedback = 32'h80000414;
            else if((index % 100) == 27) assign feedback = 32'h80000417;
            else if((index % 100) == 28) assign feedback = 32'h80000465;
            else if((index % 100) == 29) assign feedback = 32'h8000046A;
            else if((index % 100) == 30) assign feedback = 32'h80000478;
            else if((index % 100) == 31) assign feedback = 32'h800004D4;
            else if((index % 100) == 32) assign feedback = 32'h800004F3;
            else if((index % 100) == 33) assign feedback = 32'h8000050B;
            else if((index % 100) == 34) assign feedback = 32'h80000526;
            else if((index % 100) == 35) assign feedback = 32'h8000054C;
            else if((index % 100) == 36) assign feedback = 32'h800005B6;
            else if((index % 100) == 37) assign feedback = 32'h800005C1;
            else if((index % 100) == 38) assign feedback = 32'h800005EC;
            else if((index % 100) == 39) assign feedback = 32'h800005F1;
            else if((index % 100) == 40) assign feedback = 32'h8000060D;
            else if((index % 100) == 41) assign feedback = 32'h8000060E;
            else if((index % 100) == 42) assign feedback = 32'h80000629;
            else if((index % 100) == 43) assign feedback = 32'h80000638;
            else if((index % 100) == 44) assign feedback = 32'h80000662;
            else if((index % 100) == 45) assign feedback = 32'h8000066D;
            else if((index % 100) == 46) assign feedback = 32'h80000676;
            else if((index % 100) == 47) assign feedback = 32'h800006AE;
            else if((index % 100) == 48) assign feedback = 32'h800006B0;
            else if((index % 100) == 49) assign feedback = 32'h800006BC;
            else if((index % 100) == 50) assign feedback = 32'h800006D6;
            else if((index % 100) == 51) assign feedback = 32'h8000073C;
            else if((index % 100) == 52) assign feedback = 32'h80000748;
            else if((index % 100) == 53) assign feedback = 32'h80000766;
            else if((index % 100) == 54) assign feedback = 32'h8000079C;
            else if((index % 100) == 55) assign feedback = 32'h800007B7;
            else if((index % 100) == 56) assign feedback = 32'h800007C3;
            else if((index % 100) == 57) assign feedback = 32'h800007D4;
            else if((index % 100) == 58) assign feedback = 32'h800007D8;
            else if((index % 100) == 59) assign feedback = 32'h80000806;
            else if((index % 100) == 60) assign feedback = 32'h8000083F;
            else if((index % 100) == 61) assign feedback = 32'h80000850;
            else if((index % 100) == 62) assign feedback = 32'h8000088D;
            else if((index % 100) == 63) assign feedback = 32'h800008E1;
            else if((index % 100) == 64) assign feedback = 32'h80000923;
            else if((index % 100) == 65) assign feedback = 32'h80000931;
            else if((index % 100) == 66) assign feedback = 32'h80000934;
            else if((index % 100) == 67) assign feedback = 32'h8000093B;
            else if((index % 100) == 68) assign feedback = 32'h80000958;
            else if((index % 100) == 69) assign feedback = 32'h80000967;
            else if((index % 100) == 70) assign feedback = 32'h800009D5;
            else if((index % 100) == 71) assign feedback = 32'h80000A25;
            else if((index % 100) == 72) assign feedback = 32'h80000A26;
            else if((index % 100) == 73) assign feedback = 32'h80000A54;
            else if((index % 100) == 74) assign feedback = 32'h80000A92;
            else if((index % 100) == 75) assign feedback = 32'h80000AC4;
            else if((index % 100) == 76) assign feedback = 32'h80000ACD;
            else if((index % 100) == 77) assign feedback = 32'h80000B28;
            else if((index % 100) == 78) assign feedback = 32'h80000B71;
            else if((index % 100) == 79) assign feedback = 32'h80000B7B;
            else if((index % 100) == 80) assign feedback = 32'h80000B84;
            else if((index % 100) == 81) assign feedback = 32'h80000BA9;
            else if((index % 100) == 82) assign feedback = 32'h80000BBE;
            else if((index % 100) == 83) assign feedback = 32'h80000BC6;
            else if((index % 100) == 84) assign feedback = 32'h80000C34;
            else if((index % 100) == 85) assign feedback = 32'h80000C3E;
            else if((index % 100) == 86) assign feedback = 32'h80000C43;
            else if((index % 100) == 87) assign feedback = 32'h80000C7F;
            else if((index % 100) == 88) assign feedback = 32'h80000CA2;
            else if((index % 100) == 89) assign feedback = 32'h80000CEC;
            else if((index % 100) == 90) assign feedback = 32'h80000D0F;
            else if((index % 100) == 91) assign feedback = 32'h80000D22;
            else if((index % 100) == 92) assign feedback = 32'h80000D28;
            else if((index % 100) == 93) assign feedback = 32'h80000D4E;
            else if((index % 100) == 94) assign feedback = 32'h80000DD7;
            else if((index % 100) == 95) assign feedback = 32'h80000E24;
            else if((index % 100) == 96) assign feedback = 32'h80000E35;
            else if((index % 100) == 97) assign feedback = 32'h80000E66;
            else if((index % 100) == 98) assign feedback = 32'h80000E74;
            else if((index % 100) == 99) assign feedback = 32'h80000EA6;
         end
      else if(width == 33)
         begin
            if((index % 100) == 0) assign feedback = 33'h100000029;
            else if((index % 100) == 1) assign feedback = 33'h100000034;
            else if((index % 100) == 2) assign feedback = 33'h100000043;
            else if((index % 100) == 3) assign feedback = 33'h10000004C;
            else if((index % 100) == 4) assign feedback = 33'h100000051;
            else if((index % 100) == 5) assign feedback = 33'h10000006E;
            else if((index % 100) == 6) assign feedback = 33'h100000076;
            else if((index % 100) == 7) assign feedback = 33'h10000007A;
            else if((index % 100) == 8) assign feedback = 33'h100000083;
            else if((index % 100) == 9) assign feedback = 33'h100000091;
            else if((index % 100) == 10) assign feedback = 33'h100000098;
            else if((index % 100) == 11) assign feedback = 33'h1000000A7;
            else if((index % 100) == 12) assign feedback = 33'h1000000B6;
            else if((index % 100) == 13) assign feedback = 33'h1000000BC;
            else if((index % 100) == 14) assign feedback = 33'h1000000C1;
            else if((index % 100) == 15) assign feedback = 33'h1000000E3;
            else if((index % 100) == 16) assign feedback = 33'h1000000E6;
            else if((index % 100) == 17) assign feedback = 33'h1000000F1;
            else if((index % 100) == 18) assign feedback = 33'h1000000F8;
            else if((index % 100) == 19) assign feedback = 33'h1000000FE;
            else if((index % 100) == 20) assign feedback = 33'h100000105;
            else if((index % 100) == 21) assign feedback = 33'h10000010F;
            else if((index % 100) == 22) assign feedback = 33'h10000013F;
            else if((index % 100) == 23) assign feedback = 33'h10000014D;
            else if((index % 100) == 24) assign feedback = 33'h10000014E;
            else if((index % 100) == 25) assign feedback = 33'h100000153;
            else if((index % 100) == 26) assign feedback = 33'h10000015C;
            else if((index % 100) == 27) assign feedback = 33'h100000184;
            else if((index % 100) == 28) assign feedback = 33'h100000199;
            else if((index % 100) == 29) assign feedback = 33'h10000019F;
            else if((index % 100) == 30) assign feedback = 33'h1000001A3;
            else if((index % 100) == 31) assign feedback = 33'h1000001A9;
            else if((index % 100) == 32) assign feedback = 33'h1000001AF;
            else if((index % 100) == 33) assign feedback = 33'h1000001BD;
            else if((index % 100) == 34) assign feedback = 33'h1000001CC;
            else if((index % 100) == 35) assign feedback = 33'h1000001EE;
            else if((index % 100) == 36) assign feedback = 33'h1000001F5;
            else if((index % 100) == 37) assign feedback = 33'h100000203;
            else if((index % 100) == 38) assign feedback = 33'h10000021E;
            else if((index % 100) == 39) assign feedback = 33'h100000235;
            else if((index % 100) == 40) assign feedback = 33'h100000244;
            else if((index % 100) == 41) assign feedback = 33'h10000026C;
            else if((index % 100) == 42) assign feedback = 33'h100000274;
            else if((index % 100) == 43) assign feedback = 33'h10000027D;
            else if((index % 100) == 44) assign feedback = 33'h10000029A;
            else if((index % 100) == 45) assign feedback = 33'h1000002A5;
            else if((index % 100) == 46) assign feedback = 33'h1000002DB;
            else if((index % 100) == 47) assign feedback = 33'h1000002EB;
            else if((index % 100) == 48) assign feedback = 33'h10000031C;
            else if((index % 100) == 49) assign feedback = 33'h100000349;
            else if((index % 100) == 50) assign feedback = 33'h100000357;
            else if((index % 100) == 51) assign feedback = 33'h10000036B;
            else if((index % 100) == 52) assign feedback = 33'h10000036D;
            else if((index % 100) == 53) assign feedback = 33'h100000383;
            else if((index % 100) == 54) assign feedback = 33'h1000003AE;
            else if((index % 100) == 55) assign feedback = 33'h1000003EA;
            else if((index % 100) == 56) assign feedback = 33'h1000003EF;
            else if((index % 100) == 57) assign feedback = 33'h100000403;
            else if((index % 100) == 58) assign feedback = 33'h100000412;
            else if((index % 100) == 59) assign feedback = 33'h100000439;
            else if((index % 100) == 60) assign feedback = 33'h100000447;
            else if((index % 100) == 61) assign feedback = 33'h10000045A;
            else if((index % 100) == 62) assign feedback = 33'h100000478;
            else if((index % 100) == 63) assign feedback = 33'h100000484;
            else if((index % 100) == 64) assign feedback = 33'h1000004B2;
            else if((index % 100) == 65) assign feedback = 33'h1000004DB;
            else if((index % 100) == 66) assign feedback = 33'h1000004FF;
            else if((index % 100) == 67) assign feedback = 33'h100000526;
            else if((index % 100) == 68) assign feedback = 33'h10000052F;
            else if((index % 100) == 69) assign feedback = 33'h100000558;
            else if((index % 100) == 70) assign feedback = 33'h100000575;
            else if((index % 100) == 71) assign feedback = 33'h100000580;
            else if((index % 100) == 72) assign feedback = 33'h100000585;
            else if((index % 100) == 73) assign feedback = 33'h1000005A1;
            else if((index % 100) == 74) assign feedback = 33'h1000005BA;
            else if((index % 100) == 75) assign feedback = 33'h1000005DC;
            else if((index % 100) == 76) assign feedback = 33'h1000005DF;
            else if((index % 100) == 77) assign feedback = 33'h1000005F1;
            else if((index % 100) == 78) assign feedback = 33'h100000602;
            else if((index % 100) == 79) assign feedback = 33'h100000608;
            else if((index % 100) == 80) assign feedback = 33'h100000610;
            else if((index % 100) == 81) assign feedback = 33'h100000664;
            else if((index % 100) == 82) assign feedback = 33'h10000066B;
            else if((index % 100) == 83) assign feedback = 33'h100000689;
            else if((index % 100) == 84) assign feedback = 33'h1000006B3;
            else if((index % 100) == 85) assign feedback = 33'h1000006E5;
            else if((index % 100) == 86) assign feedback = 33'h1000006E6;
            else if((index % 100) == 87) assign feedback = 33'h1000006FB;
            else if((index % 100) == 88) assign feedback = 33'h100000711;
            else if((index % 100) == 89) assign feedback = 33'h100000714;
            else if((index % 100) == 90) assign feedback = 33'h100000735;
            else if((index % 100) == 91) assign feedback = 33'h10000073A;
            else if((index % 100) == 92) assign feedback = 33'h100000747;
            else if((index % 100) == 93) assign feedback = 33'h10000074B;
            else if((index % 100) == 94) assign feedback = 33'h100000763;
            else if((index % 100) == 95) assign feedback = 33'h100000766;
            else if((index % 100) == 96) assign feedback = 33'h100000769;
            else if((index % 100) == 97) assign feedback = 33'h100000784;
            else if((index % 100) == 98) assign feedback = 33'h100000788;
            else if((index % 100) == 99) assign feedback = 33'h1000007A3;
         end
      else if(width == 34)
         begin
            if((index % 100) == 0) assign feedback = 34'h200000073;
            else if((index % 100) == 1) assign feedback = 34'h20000008C;
            else if((index % 100) == 2) assign feedback = 34'h20000008F;
            else if((index % 100) == 3) assign feedback = 34'h2000000BA;
            else if((index % 100) == 4) assign feedback = 34'h2000000C7;
            else if((index % 100) == 5) assign feedback = 34'h2000000D9;
            else if((index % 100) == 6) assign feedback = 34'h2000000E9;
            else if((index % 100) == 7) assign feedback = 34'h2000000F2;
            else if((index % 100) == 8) assign feedback = 34'h200000111;
            else if((index % 100) == 9) assign feedback = 34'h200000128;
            else if((index % 100) == 10) assign feedback = 34'h20000015F;
            else if((index % 100) == 11) assign feedback = 34'h200000172;
            else if((index % 100) == 12) assign feedback = 34'h20000018E;
            else if((index % 100) == 13) assign feedback = 34'h2000001A3;
            else if((index % 100) == 14) assign feedback = 34'h2000001C6;
            else if((index % 100) == 15) assign feedback = 34'h2000001CA;
            else if((index % 100) == 16) assign feedback = 34'h2000001D4;
            else if((index % 100) == 17) assign feedback = 34'h2000001ED;
            else if((index % 100) == 18) assign feedback = 34'h200000214;
            else if((index % 100) == 19) assign feedback = 34'h200000230;
            else if((index % 100) == 20) assign feedback = 34'h20000023F;
            else if((index % 100) == 21) assign feedback = 34'h200000253;
            else if((index % 100) == 22) assign feedback = 34'h20000025A;
            else if((index % 100) == 23) assign feedback = 34'h200000284;
            else if((index % 100) == 24) assign feedback = 34'h20000028B;
            else if((index % 100) == 25) assign feedback = 34'h200000290;
            else if((index % 100) == 26) assign feedback = 34'h2000002C5;
            else if((index % 100) == 27) assign feedback = 34'h2000002D8;
            else if((index % 100) == 28) assign feedback = 34'h200000313;
            else if((index % 100) == 29) assign feedback = 34'h200000326;
            else if((index % 100) == 30) assign feedback = 34'h20000032F;
            else if((index % 100) == 31) assign feedback = 34'h200000332;
            else if((index % 100) == 32) assign feedback = 34'h200000334;
            else if((index % 100) == 33) assign feedback = 34'h20000039D;
            else if((index % 100) == 34) assign feedback = 34'h2000003B5;
            else if((index % 100) == 35) assign feedback = 34'h2000003D0;
            else if((index % 100) == 36) assign feedback = 34'h2000003DC;
            else if((index % 100) == 37) assign feedback = 34'h200000435;
            else if((index % 100) == 38) assign feedback = 34'h200000442;
            else if((index % 100) == 39) assign feedback = 34'h200000447;
            else if((index % 100) == 40) assign feedback = 34'h20000049F;
            else if((index % 100) == 41) assign feedback = 34'h2000004A5;
            else if((index % 100) == 42) assign feedback = 34'h2000004CC;
            else if((index % 100) == 43) assign feedback = 34'h200000551;
            else if((index % 100) == 44) assign feedback = 34'h20000056B;
            else if((index % 100) == 45) assign feedback = 34'h20000056E;
            else if((index % 100) == 46) assign feedback = 34'h200000575;
            else if((index % 100) == 47) assign feedback = 34'h200000580;
            else if((index % 100) == 48) assign feedback = 34'h2000005F4;
            else if((index % 100) == 49) assign feedback = 34'h2000005F7;
            else if((index % 100) == 50) assign feedback = 34'h2000005FB;
            else if((index % 100) == 51) assign feedback = 34'h2000005FE;
            else if((index % 100) == 52) assign feedback = 34'h200000626;
            else if((index % 100) == 53) assign feedback = 34'h20000062F;
            else if((index % 100) == 54) assign feedback = 34'h200000631;
            else if((index % 100) == 55) assign feedback = 34'h200000645;
            else if((index % 100) == 56) assign feedback = 34'h200000668;
            else if((index % 100) == 57) assign feedback = 34'h2000006B9;
            else if((index % 100) == 58) assign feedback = 34'h2000006D3;
            else if((index % 100) == 59) assign feedback = 34'h2000006EA;
            else if((index % 100) == 60) assign feedback = 34'h200000718;
            else if((index % 100) == 61) assign feedback = 34'h200000727;
            else if((index % 100) == 62) assign feedback = 34'h200000739;
            else if((index % 100) == 63) assign feedback = 34'h200000750;
            else if((index % 100) == 64) assign feedback = 34'h20000076A;
            else if((index % 100) == 65) assign feedback = 34'h20000076F;
            else if((index % 100) == 66) assign feedback = 34'h200000788;
            else if((index % 100) == 67) assign feedback = 34'h200000793;
            else if((index % 100) == 68) assign feedback = 34'h2000007A6;
            else if((index % 100) == 69) assign feedback = 34'h2000007C9;
            else if((index % 100) == 70) assign feedback = 34'h2000007CA;
            else if((index % 100) == 71) assign feedback = 34'h2000007ED;
            else if((index % 100) == 72) assign feedback = 34'h200000859;
            else if((index % 100) == 73) assign feedback = 34'h20000089A;
            else if((index % 100) == 74) assign feedback = 34'h2000008A6;
            else if((index % 100) == 75) assign feedback = 34'h2000008D1;
            else if((index % 100) == 76) assign feedback = 34'h2000008F0;
            else if((index % 100) == 77) assign feedback = 34'h200000904;
            else if((index % 100) == 78) assign feedback = 34'h200000925;
            else if((index % 100) == 79) assign feedback = 34'h200000929;
            else if((index % 100) == 80) assign feedback = 34'h200000932;
            else if((index % 100) == 81) assign feedback = 34'h20000093B;
            else if((index % 100) == 82) assign feedback = 34'h200000985;
            else if((index % 100) == 83) assign feedback = 34'h200000986;
            else if((index % 100) == 84) assign feedback = 34'h200000994;
            else if((index % 100) == 85) assign feedback = 34'h20000099E;
            else if((index % 100) == 86) assign feedback = 34'h2000009DC;
            else if((index % 100) == 87) assign feedback = 34'h200000A01;
            else if((index % 100) == 88) assign feedback = 34'h200000A04;
            else if((index % 100) == 89) assign feedback = 34'h200000A10;
            else if((index % 100) == 90) assign feedback = 34'h200000A26;
            else if((index % 100) == 91) assign feedback = 34'h200000A29;
            else if((index % 100) == 92) assign feedback = 34'h200000A6D;
            else if((index % 100) == 93) assign feedback = 34'h200000A73;
            else if((index % 100) == 94) assign feedback = 34'h200000A7A;
            else if((index % 100) == 95) assign feedback = 34'h200000A89;
            else if((index % 100) == 96) assign feedback = 34'h200000A94;
            else if((index % 100) == 97) assign feedback = 34'h200000AA7;
            else if((index % 100) == 98) assign feedback = 34'h200000ABC;
            else if((index % 100) == 99) assign feedback = 34'h200000ABF;
         end
      else if(width == 35)
         begin
            if((index % 93) == 0) assign feedback = 35'h400000002;
            else if((index % 93) == 1) assign feedback = 35'h40000002F;
            else if((index % 93) == 2) assign feedback = 35'h40000004F;
            else if((index % 93) == 3) assign feedback = 35'h400000057;
            else if((index % 93) == 4) assign feedback = 35'h40000009E;
            else if((index % 93) == 5) assign feedback = 35'h4000000B6;
            else if((index % 93) == 6) assign feedback = 35'h4000000C1;
            else if((index % 93) == 7) assign feedback = 35'h4000000CE;
            else if((index % 93) == 8) assign feedback = 35'h4000000DC;
            else if((index % 93) == 9) assign feedback = 35'h4000000F1;
            else if((index % 93) == 10) assign feedback = 35'h4000000F2;
            else if((index % 93) == 11) assign feedback = 35'h400000103;
            else if((index % 93) == 12) assign feedback = 35'h400000122;
            else if((index % 93) == 13) assign feedback = 35'h400000127;
            else if((index % 93) == 14) assign feedback = 35'h400000135;
            else if((index % 93) == 15) assign feedback = 35'h40000013C;
            else if((index % 93) == 16) assign feedback = 35'h400000159;
            else if((index % 93) == 17) assign feedback = 35'h400000166;
            else if((index % 93) == 18) assign feedback = 35'h400000190;
            else if((index % 93) == 19) assign feedback = 35'h4000001E4;
            else if((index % 93) == 20) assign feedback = 35'h40000020A;
            else if((index % 93) == 21) assign feedback = 35'h40000020C;
            else if((index % 93) == 22) assign feedback = 35'h400000218;
            else if((index % 93) == 23) assign feedback = 35'h400000239;
            else if((index % 93) == 24) assign feedback = 35'h400000244;
            else if((index % 93) == 25) assign feedback = 35'h40000028D;
            else if((index % 93) == 26) assign feedback = 35'h40000029A;
            else if((index % 93) == 27) assign feedback = 35'h4000002B7;
            else if((index % 93) == 28) assign feedback = 35'h4000002B8;
            else if((index % 93) == 29) assign feedback = 35'h4000002CC;
            else if((index % 93) == 30) assign feedback = 35'h4000002D2;
            else if((index % 93) == 31) assign feedback = 35'h4000002E4;
            else if((index % 93) == 32) assign feedback = 35'h4000002F0;
            else if((index % 93) == 33) assign feedback = 35'h4000002F6;
            else if((index % 93) == 34) assign feedback = 35'h4000002F9;
            else if((index % 93) == 35) assign feedback = 35'h400000301;
            else if((index % 93) == 36) assign feedback = 35'h400000308;
            else if((index % 93) == 37) assign feedback = 35'h40000032C;
            else if((index % 93) == 38) assign feedback = 35'h400000338;
            else if((index % 93) == 39) assign feedback = 35'h40000034F;
            else if((index % 93) == 40) assign feedback = 35'h40000035B;
            else if((index % 93) == 41) assign feedback = 35'h40000037F;
            else if((index % 93) == 42) assign feedback = 35'h400000380;
            else if((index % 93) == 43) assign feedback = 35'h4000003AE;
            else if((index % 93) == 44) assign feedback = 35'h4000003BA;
            else if((index % 93) == 45) assign feedback = 35'h4000003D9;
            else if((index % 93) == 46) assign feedback = 35'h400000417;
            else if((index % 93) == 47) assign feedback = 35'h40000041B;
            else if((index % 93) == 48) assign feedback = 35'h40000042D;
            else if((index % 93) == 49) assign feedback = 35'h400000430;
            else if((index % 93) == 50) assign feedback = 35'h400000453;
            else if((index % 93) == 51) assign feedback = 35'h400000463;
            else if((index % 93) == 52) assign feedback = 35'h400000471;
            else if((index % 93) == 53) assign feedback = 35'h400000478;
            else if((index % 93) == 54) assign feedback = 35'h40000048D;
            else if((index % 93) == 55) assign feedback = 35'h400000490;
            else if((index % 93) == 56) assign feedback = 35'h400000496;
            else if((index % 93) == 57) assign feedback = 35'h40000049C;
            else if((index % 93) == 58) assign feedback = 35'h4000004B2;
            else if((index % 93) == 59) assign feedback = 35'h4000004FA;
            else if((index % 93) == 60) assign feedback = 35'h40000051A;
            else if((index % 93) == 61) assign feedback = 35'h40000052C;
            else if((index % 93) == 62) assign feedback = 35'h40000055E;
            else if((index % 93) == 63) assign feedback = 35'h400000561;
            else if((index % 93) == 64) assign feedback = 35'h400000594;
            else if((index % 93) == 65) assign feedback = 35'h4000005AB;
            else if((index % 93) == 66) assign feedback = 35'h4000005AE;
            else if((index % 93) == 67) assign feedback = 35'h4000005E5;
            else if((index % 93) == 68) assign feedback = 35'h4000005E6;
            else if((index % 93) == 69) assign feedback = 35'h4000005F8;
            else if((index % 93) == 70) assign feedback = 35'h40000061F;
            else if((index % 93) == 71) assign feedback = 35'h400000623;
            else if((index % 93) == 72) assign feedback = 35'h400000631;
            else if((index % 93) == 73) assign feedback = 35'h40000063E;
            else if((index % 93) == 74) assign feedback = 35'h400000652;
            else if((index % 93) == 75) assign feedback = 35'h400000668;
            else if((index % 93) == 76) assign feedback = 35'h40000066B;
            else if((index % 93) == 77) assign feedback = 35'h400000670;
            else if((index % 93) == 78) assign feedback = 35'h4000006CE;
            else if((index % 93) == 79) assign feedback = 35'h4000006E3;
            else if((index % 93) == 80) assign feedback = 35'h400000700;
            else if((index % 93) == 81) assign feedback = 35'h400000709;
            else if((index % 93) == 82) assign feedback = 35'h400000717;
            else if((index % 93) == 83) assign feedback = 35'h40000071B;
            else if((index % 93) == 84) assign feedback = 35'h40000071E;
            else if((index % 93) == 85) assign feedback = 35'h400000728;
            else if((index % 93) == 86) assign feedback = 35'h400000777;
            else if((index % 93) == 87) assign feedback = 35'h4000007B4;
            else if((index % 93) == 88) assign feedback = 35'h4000007CF;
            else if((index % 93) == 89) assign feedback = 35'h4000007D1;
            else if((index % 93) == 90) assign feedback = 35'h4000007D2;
            else if((index % 93) == 91) assign feedback = 35'h4000007DD;
            else if((index % 93) == 92) assign feedback = 35'h4000007EB;
         end
      else if(width == 36)
         begin
            if((index % 100) == 0) assign feedback = 36'h80000003B;
            else if((index % 100) == 1) assign feedback = 36'h80000003D;
            else if((index % 100) == 2) assign feedback = 36'h80000007C;
            else if((index % 100) == 3) assign feedback = 36'h8000000B5;
            else if((index % 100) == 4) assign feedback = 36'h8000000C1;
            else if((index % 100) == 5) assign feedback = 36'h8000000F7;
            else if((index % 100) == 6) assign feedback = 36'h80000010C;
            else if((index % 100) == 7) assign feedback = 36'h80000011D;
            else if((index % 100) == 8) assign feedback = 36'h800000133;
            else if((index % 100) == 9) assign feedback = 36'h800000141;
            else if((index % 100) == 10) assign feedback = 36'h800000156;
            else if((index % 100) == 11) assign feedback = 36'h800000169;
            else if((index % 100) == 12) assign feedback = 36'h800000171;
            else if((index % 100) == 13) assign feedback = 36'h800000190;
            else if((index % 100) == 14) assign feedback = 36'h8000001B8;
            else if((index % 100) == 15) assign feedback = 36'h8000001E2;
            else if((index % 100) == 16) assign feedback = 36'h8000001FA;
            else if((index % 100) == 17) assign feedback = 36'h8000001FC;
            else if((index % 100) == 18) assign feedback = 36'h800000221;
            else if((index % 100) == 19) assign feedback = 36'h800000256;
            else if((index % 100) == 20) assign feedback = 36'h80000028B;
            else if((index % 100) == 21) assign feedback = 36'h800000299;
            else if((index % 100) == 22) assign feedback = 36'h8000002DD;
            else if((index % 100) == 23) assign feedback = 36'h80000030D;
            else if((index % 100) == 24) assign feedback = 36'h800000345;
            else if((index % 100) == 25) assign feedback = 36'h8000003A2;
            else if((index % 100) == 26) assign feedback = 36'h8000003CE;
            else if((index % 100) == 27) assign feedback = 36'h800000400;
            else if((index % 100) == 28) assign feedback = 36'h800000448;
            else if((index % 100) == 29) assign feedback = 36'h8000004CC;
            else if((index % 100) == 30) assign feedback = 36'h800000510;
            else if((index % 100) == 31) assign feedback = 36'h800000589;
            else if((index % 100) == 32) assign feedback = 36'h8000005DF;
            else if((index % 100) == 33) assign feedback = 36'h80000063D;
            else if((index % 100) == 34) assign feedback = 36'h800000667;
            else if((index % 100) == 35) assign feedback = 36'h800000676;
            else if((index % 100) == 36) assign feedback = 36'h800000697;
            else if((index % 100) == 37) assign feedback = 36'h800000772;
            else if((index % 100) == 38) assign feedback = 36'h800000778;
            else if((index % 100) == 39) assign feedback = 36'h800000787;
            else if((index % 100) == 40) assign feedback = 36'h8000007C6;
            else if((index % 100) == 41) assign feedback = 36'h800000830;
            else if((index % 100) == 42) assign feedback = 36'h800000848;
            else if((index % 100) == 43) assign feedback = 36'h800000855;
            else if((index % 100) == 44) assign feedback = 36'h80000087B;
            else if((index % 100) == 45) assign feedback = 36'h80000087E;
            else if((index % 100) == 46) assign feedback = 36'h80000088B;
            else if((index % 100) == 47) assign feedback = 36'h8000008B1;
            else if((index % 100) == 48) assign feedback = 36'h8000008BD;
            else if((index % 100) == 49) assign feedback = 36'h800000919;
            else if((index % 100) == 50) assign feedback = 36'h800000929;
            else if((index % 100) == 51) assign feedback = 36'h8000009A7;
            else if((index % 100) == 52) assign feedback = 36'h8000009DC;
            else if((index % 100) == 53) assign feedback = 36'h800000A01;
            else if((index % 100) == 54) assign feedback = 36'h800000A31;
            else if((index % 100) == 55) assign feedback = 36'h800000A32;
            else if((index % 100) == 56) assign feedback = 36'h800000A62;
            else if((index % 100) == 57) assign feedback = 36'h800000B17;
            else if((index % 100) == 58) assign feedback = 36'h800000B2E;
            else if((index % 100) == 59) assign feedback = 36'h800000B6C;
            else if((index % 100) == 60) assign feedback = 36'h800000B7E;
            else if((index % 100) == 61) assign feedback = 36'h800000B82;
            else if((index % 100) == 62) assign feedback = 36'h800000B95;
            else if((index % 100) == 63) assign feedback = 36'h800000B9A;
            else if((index % 100) == 64) assign feedback = 36'h800000B9C;
            else if((index % 100) == 65) assign feedback = 36'h800000BA6;
            else if((index % 100) == 66) assign feedback = 36'h800000BD1;
            else if((index % 100) == 67) assign feedback = 36'h800000BEB;
            else if((index % 100) == 68) assign feedback = 36'h800000C0B;
            else if((index % 100) == 69) assign feedback = 36'h800000C23;
            else if((index % 100) == 70) assign feedback = 36'h800000C51;
            else if((index % 100) == 71) assign feedback = 36'h800000C61;
            else if((index % 100) == 72) assign feedback = 36'h800000C7C;
            else if((index % 100) == 73) assign feedback = 36'h800000CCD;
            else if((index % 100) == 74) assign feedback = 36'h800000CDC;
            else if((index % 100) == 75) assign feedback = 36'h800000D65;
            else if((index % 100) == 76) assign feedback = 36'h800000D74;
            else if((index % 100) == 77) assign feedback = 36'h800000D7E;
            else if((index % 100) == 78) assign feedback = 36'h800000D99;
            else if((index % 100) == 79) assign feedback = 36'h800000DC9;
            else if((index % 100) == 80) assign feedback = 36'h800000DD8;
            else if((index % 100) == 81) assign feedback = 36'h800000E11;
            else if((index % 100) == 82) assign feedback = 36'h800000E17;
            else if((index % 100) == 83) assign feedback = 36'h800000F79;
            else if((index % 100) == 84) assign feedback = 36'h800000F89;
            else if((index % 100) == 85) assign feedback = 36'h800000F9E;
            else if((index % 100) == 86) assign feedback = 36'h800000FD9;
            else if((index % 100) == 87) assign feedback = 36'h800000FE0;
            else if((index % 100) == 88) assign feedback = 36'h800000FE6;
            else if((index % 100) == 89) assign feedback = 36'h800000FF7;
            else if((index % 100) == 90) assign feedback = 36'h800001081;
            else if((index % 100) == 91) assign feedback = 36'h8000010C0;
            else if((index % 100) == 92) assign feedback = 36'h8000010D8;
            else if((index % 100) == 93) assign feedback = 36'h80000111F;
            else if((index % 100) == 94) assign feedback = 36'h800001120;
            else if((index % 100) == 95) assign feedback = 36'h800001176;
            else if((index % 100) == 96) assign feedback = 36'h8000011D5;
            else if((index % 100) == 97) assign feedback = 36'h8000011E3;
            else if((index % 100) == 98) assign feedback = 36'h80000122F;
            else if((index % 100) == 99) assign feedback = 36'h80000123E;
         end
      else if(width == 37)
         begin
            if((index % 100) == 0) assign feedback = 37'h100000001F;
            else if((index % 100) == 1) assign feedback = 37'h1000000029;
            else if((index % 100) == 2) assign feedback = 37'h1000000038;
            else if((index % 100) == 3) assign feedback = 37'h100000005B;
            else if((index % 100) == 4) assign feedback = 37'h1000000064;
            else if((index % 100) == 5) assign feedback = 37'h1000000068;
            else if((index % 100) == 6) assign feedback = 37'h100000007A;
            else if((index % 100) == 7) assign feedback = 37'h100000009E;
            else if((index % 100) == 8) assign feedback = 37'h10000000AE;
            else if((index % 100) == 9) assign feedback = 37'h10000000C4;
            else if((index % 100) == 10) assign feedback = 37'h10000000E3;
            else if((index % 100) == 11) assign feedback = 37'h10000000E6;
            else if((index % 100) == 12) assign feedback = 37'h10000000E9;
            else if((index % 100) == 13) assign feedback = 37'h10000000F8;
            else if((index % 100) == 14) assign feedback = 37'h1000000103;
            else if((index % 100) == 15) assign feedback = 37'h100000010C;
            else if((index % 100) == 16) assign feedback = 37'h100000017D;
            else if((index % 100) == 17) assign feedback = 37'h100000019C;
            else if((index % 100) == 18) assign feedback = 37'h10000001A6;
            else if((index % 100) == 19) assign feedback = 37'h10000001AA;
            else if((index % 100) == 20) assign feedback = 37'h10000001AF;
            else if((index % 100) == 21) assign feedback = 37'h10000001B1;
            else if((index % 100) == 22) assign feedback = 37'h10000001B7;
            else if((index % 100) == 23) assign feedback = 37'h10000001CF;
            else if((index % 100) == 24) assign feedback = 37'h10000001DD;
            else if((index % 100) == 25) assign feedback = 37'h10000001F9;
            else if((index % 100) == 26) assign feedback = 37'h1000000214;
            else if((index % 100) == 27) assign feedback = 37'h1000000233;
            else if((index % 100) == 28) assign feedback = 37'h1000000260;
            else if((index % 100) == 29) assign feedback = 37'h1000000271;
            else if((index % 100) == 30) assign feedback = 37'h100000028B;
            else if((index % 100) == 31) assign feedback = 37'h100000028E;
            else if((index % 100) == 32) assign feedback = 37'h10000002B4;
            else if((index % 100) == 33) assign feedback = 37'h10000002BB;
            else if((index % 100) == 34) assign feedback = 37'h10000002DE;
            else if((index % 100) == 35) assign feedback = 37'h10000002E1;
            else if((index % 100) == 36) assign feedback = 37'h10000002E7;
            else if((index % 100) == 37) assign feedback = 37'h10000002F0;
            else if((index % 100) == 38) assign feedback = 37'h10000002F5;
            else if((index % 100) == 39) assign feedback = 37'h1000000316;
            else if((index % 100) == 40) assign feedback = 37'h1000000329;
            else if((index % 100) == 41) assign feedback = 37'h1000000332;
            else if((index % 100) == 42) assign feedback = 37'h1000000345;
            else if((index % 100) == 43) assign feedback = 37'h100000035B;
            else if((index % 100) == 44) assign feedback = 37'h100000037A;
            else if((index % 100) == 45) assign feedback = 37'h1000000386;
            else if((index % 100) == 46) assign feedback = 37'h100000038A;
            else if((index % 100) == 47) assign feedback = 37'h10000003AB;
            else if((index % 100) == 48) assign feedback = 37'h10000003B9;
            else if((index % 100) == 49) assign feedback = 37'h10000003BC;
            else if((index % 100) == 50) assign feedback = 37'h10000003D0;
            else if((index % 100) == 51) assign feedback = 37'h10000003DA;
            else if((index % 100) == 52) assign feedback = 37'h10000003EF;
            else if((index % 100) == 53) assign feedback = 37'h1000000421;
            else if((index % 100) == 54) assign feedback = 37'h1000000433;
            else if((index % 100) == 55) assign feedback = 37'h1000000442;
            else if((index % 100) == 56) assign feedback = 37'h100000044B;
            else if((index % 100) == 57) assign feedback = 37'h1000000463;
            else if((index % 100) == 58) assign feedback = 37'h1000000471;
            else if((index % 100) == 59) assign feedback = 37'h1000000472;
            else if((index % 100) == 60) assign feedback = 37'h100000049C;
            else if((index % 100) == 61) assign feedback = 37'h10000004AC;
            else if((index % 100) == 62) assign feedback = 37'h10000004B1;
            else if((index % 100) == 63) assign feedback = 37'h10000004BE;
            else if((index % 100) == 64) assign feedback = 37'h10000004C9;
            else if((index % 100) == 65) assign feedback = 37'h10000004D7;
            else if((index % 100) == 66) assign feedback = 37'h10000004E1;
            else if((index % 100) == 67) assign feedback = 37'h10000004E4;
            else if((index % 100) == 68) assign feedback = 37'h10000004F6;
            else if((index % 100) == 69) assign feedback = 37'h10000004F9;
            else if((index % 100) == 70) assign feedback = 37'h1000000523;
            else if((index % 100) == 71) assign feedback = 37'h1000000526;
            else if((index % 100) == 72) assign feedback = 37'h100000054F;
            else if((index % 100) == 73) assign feedback = 37'h1000000562;
            else if((index % 100) == 74) assign feedback = 37'h1000000575;
            else if((index % 100) == 75) assign feedback = 37'h1000000592;
            else if((index % 100) == 76) assign feedback = 37'h10000005BC;
            else if((index % 100) == 77) assign feedback = 37'h10000005C1;
            else if((index % 100) == 78) assign feedback = 37'h10000005C8;
            else if((index % 100) == 79) assign feedback = 37'h10000005DA;
            else if((index % 100) == 80) assign feedback = 37'h10000005E0;
            else if((index % 100) == 81) assign feedback = 37'h10000005F4;
            else if((index % 100) == 82) assign feedback = 37'h100000060D;
            else if((index % 100) == 83) assign feedback = 37'h1000000623;
            else if((index % 100) == 84) assign feedback = 37'h1000000632;
            else if((index % 100) == 85) assign feedback = 37'h1000000634;
            else if((index % 100) == 86) assign feedback = 37'h100000066B;
            else if((index % 100) == 87) assign feedback = 37'h100000066E;
            else if((index % 100) == 88) assign feedback = 37'h1000000679;
            else if((index % 100) == 89) assign feedback = 37'h1000000680;
            else if((index % 100) == 90) assign feedback = 37'h100000069B;
            else if((index % 100) == 91) assign feedback = 37'h10000006A1;
            else if((index % 100) == 92) assign feedback = 37'h10000006AB;
            else if((index % 100) == 93) assign feedback = 37'h10000006D6;
            else if((index % 100) == 94) assign feedback = 37'h10000006DF;
            else if((index % 100) == 95) assign feedback = 37'h10000006F1;
            else if((index % 100) == 96) assign feedback = 37'h10000006F2;
            else if((index % 100) == 97) assign feedback = 37'h1000000718;
            else if((index % 100) == 98) assign feedback = 37'h1000000722;
            else if((index % 100) == 99) assign feedback = 37'h100000074E;
         end
      else if(width == 38)
         begin
            if((index % 100) == 0) assign feedback = 38'h2000000031;
            else if((index % 100) == 1) assign feedback = 38'h2000000051;
            else if((index % 100) == 2) assign feedback = 38'h200000006B;
            else if((index % 100) == 3) assign feedback = 38'h20000000A1;
            else if((index % 100) == 4) assign feedback = 38'h20000000B9;
            else if((index % 100) == 5) assign feedback = 38'h20000000D5;
            else if((index % 100) == 6) assign feedback = 38'h20000000F8;
            else if((index % 100) == 7) assign feedback = 38'h20000000FB;
            else if((index % 100) == 8) assign feedback = 38'h2000000106;
            else if((index % 100) == 9) assign feedback = 38'h2000000163;
            else if((index % 100) == 10) assign feedback = 38'h2000000184;
            else if((index % 100) == 11) assign feedback = 38'h2000000199;
            else if((index % 100) == 12) assign feedback = 38'h20000001B2;
            else if((index % 100) == 13) assign feedback = 38'h20000001B4;
            else if((index % 100) == 14) assign feedback = 38'h200000020F;
            else if((index % 100) == 15) assign feedback = 38'h2000000239;
            else if((index % 100) == 16) assign feedback = 38'h200000026F;
            else if((index % 100) == 17) assign feedback = 38'h200000027D;
            else if((index % 100) == 18) assign feedback = 38'h20000002AC;
            else if((index % 100) == 19) assign feedback = 38'h20000002B2;
            else if((index % 100) == 20) assign feedback = 38'h20000002B8;
            else if((index % 100) == 21) assign feedback = 38'h200000032F;
            else if((index % 100) == 22) assign feedback = 38'h2000000334;
            else if((index % 100) == 23) assign feedback = 38'h200000037C;
            else if((index % 100) == 24) assign feedback = 38'h200000037F;
            else if((index % 100) == 25) assign feedback = 38'h2000000389;
            else if((index % 100) == 26) assign feedback = 38'h2000000398;
            else if((index % 100) == 27) assign feedback = 38'h20000003A8;
            else if((index % 100) == 28) assign feedback = 38'h20000003C1;
            else if((index % 100) == 29) assign feedback = 38'h20000003CB;
            else if((index % 100) == 30) assign feedback = 38'h20000003CD;
            else if((index % 100) == 31) assign feedback = 38'h20000003DA;
            else if((index % 100) == 32) assign feedback = 38'h2000000412;
            else if((index % 100) == 33) assign feedback = 38'h200000041B;
            else if((index % 100) == 34) assign feedback = 38'h2000000428;
            else if((index % 100) == 35) assign feedback = 38'h200000043F;
            else if((index % 100) == 36) assign feedback = 38'h200000046A;
            else if((index % 100) == 37) assign feedback = 38'h2000000472;
            else if((index % 100) == 38) assign feedback = 38'h2000000477;
            else if((index % 100) == 39) assign feedback = 38'h2000000490;
            else if((index % 100) == 40) assign feedback = 38'h20000004AA;
            else if((index % 100) == 41) assign feedback = 38'h20000004BD;
            else if((index % 100) == 42) assign feedback = 38'h20000004C5;
            else if((index % 100) == 43) assign feedback = 38'h20000004DE;
            else if((index % 100) == 44) assign feedback = 38'h200000051A;
            else if((index % 100) == 45) assign feedback = 38'h2000000552;
            else if((index % 100) == 46) assign feedback = 38'h200000055B;
            else if((index % 100) == 47) assign feedback = 38'h2000000564;
            else if((index % 100) == 48) assign feedback = 38'h2000000568;
            else if((index % 100) == 49) assign feedback = 38'h2000000573;
            else if((index % 100) == 50) assign feedback = 38'h20000005D3;
            else if((index % 100) == 51) assign feedback = 38'h20000005DC;
            else if((index % 100) == 52) assign feedback = 38'h20000005E6;
            else if((index % 100) == 53) assign feedback = 38'h20000005EF;
            else if((index % 100) == 54) assign feedback = 38'h20000005FD;
            else if((index % 100) == 55) assign feedback = 38'h2000000640;
            else if((index % 100) == 56) assign feedback = 38'h2000000646;
            else if((index % 100) == 57) assign feedback = 38'h200000064F;
            else if((index % 100) == 58) assign feedback = 38'h2000000657;
            else if((index % 100) == 59) assign feedback = 38'h2000000694;
            else if((index % 100) == 60) assign feedback = 38'h2000000709;
            else if((index % 100) == 61) assign feedback = 38'h2000000711;
            else if((index % 100) == 62) assign feedback = 38'h200000072D;
            else if((index % 100) == 63) assign feedback = 38'h2000000742;
            else if((index % 100) == 64) assign feedback = 38'h2000000756;
            else if((index % 100) == 65) assign feedback = 38'h200000076F;
            else if((index % 100) == 66) assign feedback = 38'h200000078B;
            else if((index % 100) == 67) assign feedback = 38'h2000000795;
            else if((index % 100) == 68) assign feedback = 38'h20000007AC;
            else if((index % 100) == 69) assign feedback = 38'h20000007B8;
            else if((index % 100) == 70) assign feedback = 38'h20000007BE;
            else if((index % 100) == 71) assign feedback = 38'h20000007E2;
            else if((index % 100) == 72) assign feedback = 38'h20000007EE;
            else if((index % 100) == 73) assign feedback = 38'h20000007FC;
            else if((index % 100) == 74) assign feedback = 38'h2000000818;
            else if((index % 100) == 75) assign feedback = 38'h200000081B;
            else if((index % 100) == 76) assign feedback = 38'h200000081D;
            else if((index % 100) == 77) assign feedback = 38'h200000083F;
            else if((index % 100) == 78) assign feedback = 38'h200000085C;
            else if((index % 100) == 79) assign feedback = 38'h20000008AF;
            else if((index % 100) == 80) assign feedback = 38'h20000008B4;
            else if((index % 100) == 81) assign feedback = 38'h2000000902;
            else if((index % 100) == 82) assign feedback = 38'h200000090D;
            else if((index % 100) == 83) assign feedback = 38'h200000091C;
            else if((index % 100) == 84) assign feedback = 38'h2000000926;
            else if((index % 100) == 85) assign feedback = 38'h2000000980;
            else if((index % 100) == 86) assign feedback = 38'h2000000989;
            else if((index % 100) == 87) assign feedback = 38'h20000009A1;
            else if((index % 100) == 88) assign feedback = 38'h20000009AD;
            else if((index % 100) == 89) assign feedback = 38'h20000009BA;
            else if((index % 100) == 90) assign feedback = 38'h20000009C8;
            else if((index % 100) == 91) assign feedback = 38'h2000000A37;
            else if((index % 100) == 92) assign feedback = 38'h2000000A54;
            else if((index % 100) == 93) assign feedback = 38'h2000000A6D;
            else if((index % 100) == 94) assign feedback = 38'h2000000A6E;
            else if((index % 100) == 95) assign feedback = 38'h2000000AA4;
            else if((index % 100) == 96) assign feedback = 38'h2000000AC4;
            else if((index % 100) == 97) assign feedback = 38'h2000000AC8;
            else if((index % 100) == 98) assign feedback = 38'h2000000ACD;
            else if((index % 100) == 99) assign feedback = 38'h2000000AE9;
         end
      else if(width == 39)
         begin
            if((index % 61) == 0) assign feedback = 39'h4000000008;
            else if((index % 61) == 1) assign feedback = 39'h4000000049;
            else if((index % 61) == 2) assign feedback = 39'h400000006E;
            else if((index % 61) == 3) assign feedback = 39'h4000000080;
            else if((index % 61) == 4) assign feedback = 39'h40000000A4;
            else if((index % 61) == 5) assign feedback = 39'h40000000E3;
            else if((index % 61) == 6) assign feedback = 39'h40000000F1;
            else if((index % 61) == 7) assign feedback = 39'h4000000105;
            else if((index % 61) == 8) assign feedback = 39'h4000000106;
            else if((index % 61) == 9) assign feedback = 39'h4000000117;
            else if((index % 61) == 10) assign feedback = 39'h4000000121;
            else if((index % 61) == 11) assign feedback = 39'h400000012D;
            else if((index % 61) == 12) assign feedback = 39'h4000000130;
            else if((index % 61) == 13) assign feedback = 39'h400000013A;
            else if((index % 61) == 14) assign feedback = 39'h400000013F;
            else if((index % 61) == 15) assign feedback = 39'h400000014E;
            else if((index % 61) == 16) assign feedback = 39'h4000000155;
            else if((index % 61) == 17) assign feedback = 39'h4000000160;
            else if((index % 61) == 18) assign feedback = 39'h4000000172;
            else if((index % 61) == 19) assign feedback = 39'h4000000199;
            else if((index % 61) == 20) assign feedback = 39'h40000001BB;
            else if((index % 61) == 21) assign feedback = 39'h40000001CC;
            else if((index % 61) == 22) assign feedback = 39'h40000001F9;
            else if((index % 61) == 23) assign feedback = 39'h4000000227;
            else if((index % 61) == 24) assign feedback = 39'h4000000277;
            else if((index % 61) == 25) assign feedback = 39'h40000002A3;
            else if((index % 61) == 26) assign feedback = 39'h40000002AC;
            else if((index % 61) == 27) assign feedback = 39'h40000002C9;
            else if((index % 61) == 28) assign feedback = 39'h40000002D8;
            else if((index % 61) == 29) assign feedback = 39'h40000002DD;
            else if((index % 61) == 30) assign feedback = 39'h40000002F6;
            else if((index % 61) == 31) assign feedback = 39'h4000000313;
            else if((index % 61) == 32) assign feedback = 39'h400000031A;
            else if((index % 61) == 33) assign feedback = 39'h400000031C;
            else if((index % 61) == 34) assign feedback = 39'h4000000323;
            else if((index % 61) == 35) assign feedback = 39'h4000000338;
            else if((index % 61) == 36) assign feedback = 39'h4000000357;
            else if((index % 61) == 37) assign feedback = 39'h4000000361;
            else if((index % 61) == 38) assign feedback = 39'h4000000368;
            else if((index % 61) == 39) assign feedback = 39'h4000000383;
            else if((index % 61) == 40) assign feedback = 39'h4000000391;
            else if((index % 61) == 41) assign feedback = 39'h400000039D;
            else if((index % 61) == 42) assign feedback = 39'h40000003B5;
            else if((index % 61) == 43) assign feedback = 39'h40000003CE;
            else if((index % 61) == 44) assign feedback = 39'h40000003D0;
            else if((index % 61) == 45) assign feedback = 39'h40000003EF;
            else if((index % 61) == 46) assign feedback = 39'h40000003F2;
            else if((index % 61) == 47) assign feedback = 39'h400000042E;
            else if((index % 61) == 48) assign feedback = 39'h4000000441;
            else if((index % 61) == 49) assign feedback = 39'h4000000459;
            else if((index % 61) == 50) assign feedback = 39'h400000046A;
            else if((index % 61) == 51) assign feedback = 39'h400000048B;
            else if((index % 61) == 52) assign feedback = 39'h40000004A5;
            else if((index % 61) == 53) assign feedback = 39'h40000004D2;
            else if((index % 61) == 54) assign feedback = 39'h40000004E4;
            else if((index % 61) == 55) assign feedback = 39'h40000004E8;
            else if((index % 61) == 56) assign feedback = 39'h40000004F6;
            else if((index % 61) == 57) assign feedback = 39'h4000000502;
            else if((index % 61) == 58) assign feedback = 39'h400000050D;
            else if((index % 61) == 59) assign feedback = 39'h400000051C;
            else if((index % 61) == 60) assign feedback = 39'h4000000523;
         end
      // synopsys translate_off
      else
        begin
          initial
            begin
              $display("ERROR: LFSR feedback generator module %m does not support width %d.", width);
              $stop;
            end
        end
      // synopsys translate_on
      
   endgenerate
   
endmodule
